* Netlist to evaluate MOS ID-VDS characteristics
.include TSMC_180nm.txt
.param LAMBDA=0.09u
.param width_N={20*LAMBDA}

.global gnd

VGS G gnd 1.8V
VDS D gnd 0V

* MOS transistor
M1 D G gnd gnd CMOSN W={width_N} L={4*LAMBDA} 
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
+ AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

.dc VDS 0 1.8 0.1

.control
run

let id = -i(VDS)
plot id vs v(D)
.endc