.include TSMC_180nm.txt
.param Wn=1.8u
.param Wp={2.5*Wn}
.param L=0.18u
.subckt inverter in out vdd gnd Wn={Wn} Wp={Wp} L={L}
M1 out in gnd gnd CMOSN W={Wn} L={L}
M2 out in vdd vdd CMOSP W={Wp} L={L}
.ends inverter
Vdd vdd 0 1.8
Vin A 0 PWL(0n 0V 0.5n 1.8V 1.1n 1.8V 1.5n 0V 5n 0V)
Xinv1 A B vdd 0 inverter Wn={Wn} Wp={Wp} L={L}
.param scale=1
Xinv2 B C vdd 0 inverter Wn={scale*Wn} Wp={scale*Wp} L={L}
.control
tran 10p 5n
meas tran tplh TRIG v(A) VAL=0.9 RISE=1 TARG v(B) VAL=0.9 RISE=1
meas tran tphl TRIG v(A) VAL=0.9 FALL=1 TARG v(B) VAL=0.9 FALL=1
let tpd =(tplh + tphl)/2
print tpd
.endc
.end