magic
tech scmos
timestamp 1757597755
<< nwell >>
rect -14 -10 17 36
rect 24 -10 55 36
rect 62 -10 93 36
rect 100 -10 131 36
rect 138 -10 169 36
rect 176 -10 207 36
rect 214 -10 245 36
rect 252 -10 283 36
rect 290 -10 321 36
rect 328 -10 359 36
rect 366 -10 397 36
rect 404 -10 435 36
rect 442 -10 473 36
rect 480 -10 511 36
rect 518 -10 549 36
rect 556 -10 587 36
rect 594 -10 625 36
rect 632 -10 663 36
rect 670 -10 701 36
rect 708 -10 739 36
rect 746 -10 777 36
rect 784 -10 815 36
rect 822 -10 853 36
rect 860 -10 891 36
rect 898 -10 929 36
rect 936 -10 967 36
rect 974 -10 1005 36
rect 1012 -10 1043 36
rect 1050 -10 1081 36
rect 1088 -10 1119 36
rect 1126 -10 1157 36
<< ntransistor >>
rect 0 -27 2 -17
rect 38 -27 40 -17
rect 76 -27 78 -17
rect 114 -27 116 -17
rect 152 -27 154 -17
rect 190 -27 192 -17
rect 228 -27 230 -17
rect 266 -27 268 -17
rect 304 -27 306 -17
rect 342 -27 344 -17
rect 380 -27 382 -17
rect 418 -27 420 -17
rect 456 -27 458 -17
rect 494 -27 496 -17
rect 532 -27 534 -17
rect 570 -27 572 -17
rect 608 -27 610 -17
rect 646 -27 648 -17
rect 684 -27 686 -17
rect 722 -27 724 -17
rect 760 -27 762 -17
rect 798 -27 800 -17
rect 836 -27 838 -17
rect 874 -27 876 -17
rect 912 -27 914 -17
rect 950 -27 952 -17
rect 988 -27 990 -17
rect 1026 -27 1028 -17
rect 1064 -27 1066 -17
rect 1102 -27 1104 -17
rect 1140 -27 1142 -17
<< ptransistor >>
rect 0 1 2 26
rect 38 1 40 26
rect 76 1 78 26
rect 114 1 116 26
rect 152 1 154 26
rect 190 1 192 26
rect 228 1 230 26
rect 266 1 268 26
rect 304 1 306 26
rect 342 1 344 26
rect 380 1 382 26
rect 418 1 420 26
rect 456 1 458 26
rect 494 1 496 26
rect 532 1 534 26
rect 570 1 572 26
rect 608 1 610 26
rect 646 1 648 26
rect 684 1 686 26
rect 722 1 724 26
rect 760 1 762 26
rect 798 1 800 26
rect 836 1 838 26
rect 874 1 876 26
rect 912 1 914 26
rect 950 1 952 26
rect 988 1 990 26
rect 1026 1 1028 26
rect 1064 1 1066 26
rect 1102 1 1104 26
rect 1140 1 1142 26
<< ndiffusion >>
rect -3 -27 0 -17
rect 2 -27 6 -17
rect 35 -27 38 -17
rect 40 -27 44 -17
rect 73 -27 76 -17
rect 78 -27 82 -17
rect 111 -27 114 -17
rect 116 -27 120 -17
rect 149 -27 152 -17
rect 154 -27 158 -17
rect 187 -27 190 -17
rect 192 -27 196 -17
rect 225 -27 228 -17
rect 230 -27 234 -17
rect 263 -27 266 -17
rect 268 -27 272 -17
rect 301 -27 304 -17
rect 306 -27 310 -17
rect 339 -27 342 -17
rect 344 -27 348 -17
rect 377 -27 380 -17
rect 382 -27 386 -17
rect 415 -27 418 -17
rect 420 -27 424 -17
rect 453 -27 456 -17
rect 458 -27 462 -17
rect 491 -27 494 -17
rect 496 -27 500 -17
rect 529 -27 532 -17
rect 534 -27 538 -17
rect 567 -27 570 -17
rect 572 -27 576 -17
rect 605 -27 608 -17
rect 610 -27 614 -17
rect 643 -27 646 -17
rect 648 -27 652 -17
rect 681 -27 684 -17
rect 686 -27 690 -17
rect 719 -27 722 -17
rect 724 -27 728 -17
rect 757 -27 760 -17
rect 762 -27 766 -17
rect 795 -27 798 -17
rect 800 -27 804 -17
rect 833 -27 836 -17
rect 838 -27 842 -17
rect 871 -27 874 -17
rect 876 -27 880 -17
rect 909 -27 912 -17
rect 914 -27 918 -17
rect 947 -27 950 -17
rect 952 -27 956 -17
rect 985 -27 988 -17
rect 990 -27 994 -17
rect 1023 -27 1026 -17
rect 1028 -27 1032 -17
rect 1061 -27 1064 -17
rect 1066 -27 1070 -17
rect 1099 -27 1102 -17
rect 1104 -27 1108 -17
rect 1137 -27 1140 -17
rect 1142 -27 1146 -17
<< pdiffusion >>
rect -3 1 0 26
rect 2 1 6 26
rect 35 1 38 26
rect 40 1 44 26
rect 73 1 76 26
rect 78 1 82 26
rect 111 1 114 26
rect 116 1 120 26
rect 149 1 152 26
rect 154 1 158 26
rect 187 1 190 26
rect 192 1 196 26
rect 225 1 228 26
rect 230 1 234 26
rect 263 1 266 26
rect 268 1 272 26
rect 301 1 304 26
rect 306 1 310 26
rect 339 1 342 26
rect 344 1 348 26
rect 377 1 380 26
rect 382 1 386 26
rect 415 1 418 26
rect 420 1 424 26
rect 453 1 456 26
rect 458 1 462 26
rect 491 1 494 26
rect 496 1 500 26
rect 529 1 532 26
rect 534 1 538 26
rect 567 1 570 26
rect 572 1 576 26
rect 605 1 608 26
rect 610 1 614 26
rect 643 1 646 26
rect 648 1 652 26
rect 681 1 684 26
rect 686 1 690 26
rect 719 1 722 26
rect 724 1 728 26
rect 757 1 760 26
rect 762 1 766 26
rect 795 1 798 26
rect 800 1 804 26
rect 833 1 836 26
rect 838 1 842 26
rect 871 1 874 26
rect 876 1 880 26
rect 909 1 912 26
rect 914 1 918 26
rect 947 1 950 26
rect 952 1 956 26
rect 985 1 988 26
rect 990 1 994 26
rect 1023 1 1026 26
rect 1028 1 1032 26
rect 1061 1 1064 26
rect 1066 1 1070 26
rect 1099 1 1102 26
rect 1104 1 1108 26
rect 1137 1 1140 26
rect 1142 1 1146 26
<< ndcontact >>
rect -7 -27 -3 -17
rect 6 -27 10 -17
rect 31 -27 35 -17
rect 44 -27 48 -17
rect 69 -27 73 -17
rect 82 -27 86 -17
rect 107 -27 111 -17
rect 120 -27 124 -17
rect 145 -27 149 -17
rect 158 -27 162 -17
rect 183 -27 187 -17
rect 196 -27 200 -17
rect 221 -27 225 -17
rect 234 -27 238 -17
rect 259 -27 263 -17
rect 272 -27 276 -17
rect 297 -27 301 -17
rect 310 -27 314 -17
rect 335 -27 339 -17
rect 348 -27 352 -17
rect 373 -27 377 -17
rect 386 -27 390 -17
rect 411 -27 415 -17
rect 424 -27 428 -17
rect 449 -27 453 -17
rect 462 -27 466 -17
rect 487 -27 491 -17
rect 500 -27 504 -17
rect 525 -27 529 -17
rect 538 -27 542 -17
rect 563 -27 567 -17
rect 576 -27 580 -17
rect 601 -27 605 -17
rect 614 -27 618 -17
rect 639 -27 643 -17
rect 652 -27 656 -17
rect 677 -27 681 -17
rect 690 -27 694 -17
rect 715 -27 719 -17
rect 728 -27 732 -17
rect 753 -27 757 -17
rect 766 -27 770 -17
rect 791 -27 795 -17
rect 804 -27 808 -17
rect 829 -27 833 -17
rect 842 -27 846 -17
rect 867 -27 871 -17
rect 880 -27 884 -17
rect 905 -27 909 -17
rect 918 -27 922 -17
rect 943 -27 947 -17
rect 956 -27 960 -17
rect 981 -27 985 -17
rect 994 -27 998 -17
rect 1019 -27 1023 -17
rect 1032 -27 1036 -17
rect 1057 -27 1061 -17
rect 1070 -27 1074 -17
rect 1095 -27 1099 -17
rect 1108 -27 1112 -17
rect 1133 -27 1137 -17
rect 1146 -27 1150 -17
<< pdcontact >>
rect -7 1 -3 26
rect 6 1 10 26
rect 31 1 35 26
rect 44 1 48 26
rect 69 1 73 26
rect 82 1 86 26
rect 107 1 111 26
rect 120 1 124 26
rect 145 1 149 26
rect 158 1 162 26
rect 183 1 187 26
rect 196 1 200 26
rect 221 1 225 26
rect 234 1 238 26
rect 259 1 263 26
rect 272 1 276 26
rect 297 1 301 26
rect 310 1 314 26
rect 335 1 339 26
rect 348 1 352 26
rect 373 1 377 26
rect 386 1 390 26
rect 411 1 415 26
rect 424 1 428 26
rect 449 1 453 26
rect 462 1 466 26
rect 487 1 491 26
rect 500 1 504 26
rect 525 1 529 26
rect 538 1 542 26
rect 563 1 567 26
rect 576 1 580 26
rect 601 1 605 26
rect 614 1 618 26
rect 639 1 643 26
rect 652 1 656 26
rect 677 1 681 26
rect 690 1 694 26
rect 715 1 719 26
rect 728 1 732 26
rect 753 1 757 26
rect 766 1 770 26
rect 791 1 795 26
rect 804 1 808 26
rect 829 1 833 26
rect 842 1 846 26
rect 867 1 871 26
rect 880 1 884 26
rect 905 1 909 26
rect 918 1 922 26
rect 943 1 947 26
rect 956 1 960 26
rect 981 1 985 26
rect 994 1 998 26
rect 1019 1 1023 26
rect 1032 1 1036 26
rect 1057 1 1061 26
rect 1070 1 1074 26
rect 1095 1 1099 26
rect 1108 1 1112 26
rect 1133 1 1137 26
rect 1146 1 1150 26
<< polysilicon >>
rect 0 26 2 30
rect 38 26 40 30
rect 76 26 78 30
rect 114 26 116 30
rect 152 26 154 30
rect 190 26 192 30
rect 228 26 230 30
rect 266 26 268 30
rect 304 26 306 30
rect 342 26 344 30
rect 380 26 382 30
rect 418 26 420 30
rect 456 26 458 30
rect 494 26 496 30
rect 532 26 534 30
rect 570 26 572 30
rect 608 26 610 30
rect 646 26 648 30
rect 684 26 686 30
rect 722 26 724 30
rect 760 26 762 30
rect 798 26 800 30
rect 836 26 838 30
rect 874 26 876 30
rect 912 26 914 30
rect 950 26 952 30
rect 988 26 990 30
rect 1026 26 1028 30
rect 1064 26 1066 30
rect 1102 26 1104 30
rect 1140 26 1142 30
rect 0 -17 2 1
rect 38 -17 40 1
rect 76 -17 78 1
rect 114 -17 116 1
rect 152 -17 154 1
rect 190 -17 192 1
rect 228 -17 230 1
rect 266 -17 268 1
rect 304 -17 306 1
rect 342 -17 344 1
rect 380 -17 382 1
rect 418 -17 420 1
rect 456 -17 458 1
rect 494 -17 496 1
rect 532 -17 534 1
rect 570 -17 572 1
rect 608 -17 610 1
rect 646 -17 648 1
rect 684 -17 686 1
rect 722 -17 724 1
rect 760 -17 762 1
rect 798 -17 800 1
rect 836 -17 838 1
rect 874 -17 876 1
rect 912 -17 914 1
rect 950 -17 952 1
rect 988 -17 990 1
rect 1026 -17 1028 1
rect 1064 -17 1066 1
rect 1102 -17 1104 1
rect 1140 -17 1142 1
rect 0 -35 2 -27
rect 38 -35 40 -27
rect 76 -35 78 -27
rect 114 -35 116 -27
rect 152 -35 154 -27
rect 190 -35 192 -27
rect 228 -35 230 -27
rect 266 -35 268 -27
rect 304 -35 306 -27
rect 342 -35 344 -27
rect 380 -35 382 -27
rect 418 -35 420 -27
rect 456 -35 458 -27
rect 494 -35 496 -27
rect 532 -35 534 -27
rect 570 -35 572 -27
rect 608 -35 610 -27
rect 646 -35 648 -27
rect 684 -35 686 -27
rect 722 -35 724 -27
rect 760 -35 762 -27
rect 798 -35 800 -27
rect 836 -35 838 -27
rect 874 -35 876 -27
rect 912 -35 914 -27
rect 950 -35 952 -27
rect 988 -35 990 -27
rect 1026 -35 1028 -27
rect 1064 -35 1066 -27
rect 1102 -35 1104 -27
rect 1140 -35 1142 -27
<< polycontact >>
rect -4 -14 0 -10
rect 34 -14 38 -10
rect 72 -14 76 -10
rect 110 -14 114 -10
rect 148 -14 152 -10
rect 186 -14 190 -10
rect 224 -14 228 -10
rect 262 -14 266 -10
rect 300 -14 304 -10
rect 338 -14 342 -10
rect 376 -14 380 -10
rect 414 -14 418 -10
rect 452 -14 456 -10
rect 490 -14 494 -10
rect 528 -14 532 -10
rect 566 -14 570 -10
rect 604 -14 608 -10
rect 642 -14 646 -10
rect 680 -14 684 -10
rect 718 -14 722 -10
rect 756 -14 760 -10
rect 794 -14 798 -10
rect 832 -14 836 -10
rect 870 -14 874 -10
rect 908 -14 912 -10
rect 946 -14 950 -10
rect 984 -14 988 -10
rect 1022 -14 1026 -10
rect 1060 -14 1064 -10
rect 1098 -14 1102 -10
rect 1136 -14 1140 -10
<< metal1 >>
rect -28 42 1173 46
rect -28 -10 -24 42
rect -17 35 1161 39
rect -7 26 -3 35
rect 31 26 35 35
rect 69 26 73 35
rect 107 26 111 35
rect 145 26 149 35
rect 183 26 187 35
rect 221 26 225 35
rect 259 26 263 35
rect 297 26 301 35
rect 335 26 339 35
rect 373 26 377 35
rect 411 26 415 35
rect 449 26 453 35
rect 487 26 491 35
rect 525 26 529 35
rect 563 26 567 35
rect 601 26 605 35
rect 639 26 643 35
rect 677 26 681 35
rect 715 26 719 35
rect 753 26 757 35
rect 791 26 795 35
rect 829 26 833 35
rect 867 26 871 35
rect 905 26 909 35
rect 943 26 947 35
rect 981 26 985 35
rect 1019 26 1023 35
rect 1057 26 1061 35
rect 1095 26 1099 35
rect 1133 26 1137 35
rect 6 -10 10 1
rect 44 -10 48 1
rect 82 -10 86 1
rect 120 -10 124 1
rect 158 -10 162 1
rect 196 -10 200 1
rect 234 -10 238 1
rect 272 -10 276 1
rect 310 -10 314 1
rect 348 -10 352 1
rect 386 -10 390 1
rect 424 -10 428 1
rect 462 -10 466 1
rect 500 -10 504 1
rect 538 -10 542 1
rect 576 -10 580 1
rect 614 -10 618 1
rect 652 -10 656 1
rect 690 -10 694 1
rect 728 -10 732 1
rect 766 -10 770 1
rect 804 -10 808 1
rect 842 -10 846 1
rect 880 -10 884 1
rect 918 -10 922 1
rect 956 -10 960 1
rect 994 -10 998 1
rect 1032 -10 1036 1
rect 1070 -10 1074 1
rect 1108 -10 1112 1
rect 1146 -10 1150 1
rect 1168 -10 1173 42
rect -28 -14 -4 -10
rect 6 -14 34 -10
rect 44 -14 72 -10
rect 82 -14 110 -10
rect 120 -14 148 -10
rect 158 -14 186 -10
rect 196 -14 224 -10
rect 234 -14 262 -10
rect 272 -14 300 -10
rect 310 -14 338 -10
rect 348 -14 376 -10
rect 386 -14 414 -10
rect 424 -14 452 -10
rect 462 -14 490 -10
rect 500 -14 528 -10
rect 538 -14 566 -10
rect 576 -14 604 -10
rect 614 -14 642 -10
rect 652 -14 680 -10
rect 690 -14 718 -10
rect 728 -14 756 -10
rect 766 -14 794 -10
rect 804 -14 832 -10
rect 842 -14 870 -10
rect 880 -14 908 -10
rect 918 -14 946 -10
rect 956 -14 984 -10
rect 994 -14 1022 -10
rect 1032 -14 1060 -10
rect 1070 -14 1098 -10
rect 1108 -14 1136 -10
rect 1146 -14 1173 -10
rect 6 -17 10 -14
rect 44 -17 48 -14
rect 82 -17 86 -14
rect 120 -17 124 -14
rect 158 -17 162 -14
rect 196 -17 200 -14
rect 234 -17 238 -14
rect 272 -17 276 -14
rect 310 -17 314 -14
rect 348 -17 352 -14
rect 386 -17 390 -14
rect 424 -17 428 -14
rect 462 -17 466 -14
rect 500 -17 504 -14
rect 538 -17 542 -14
rect 576 -17 580 -14
rect 614 -17 618 -14
rect 652 -17 656 -14
rect 690 -17 694 -14
rect 728 -17 732 -14
rect 766 -17 770 -14
rect 804 -17 808 -14
rect 842 -17 846 -14
rect 880 -17 884 -14
rect 918 -17 922 -14
rect 956 -17 960 -14
rect 994 -17 998 -14
rect 1032 -17 1036 -14
rect 1070 -17 1074 -14
rect 1108 -17 1112 -14
rect 1146 -17 1150 -14
rect -7 -40 -3 -27
rect 31 -40 35 -27
rect 69 -40 73 -27
rect 107 -40 111 -27
rect 145 -40 149 -27
rect 183 -40 187 -27
rect 221 -40 225 -27
rect 259 -40 263 -27
rect 297 -40 301 -27
rect 335 -40 339 -27
rect 373 -40 377 -27
rect 411 -40 415 -27
rect 449 -40 453 -27
rect 487 -40 491 -27
rect 525 -40 529 -27
rect 563 -40 567 -27
rect 601 -40 605 -27
rect 639 -40 643 -27
rect 677 -40 681 -27
rect 715 -40 719 -27
rect 753 -40 757 -27
rect 791 -40 795 -27
rect 829 -40 833 -27
rect 867 -40 871 -27
rect 905 -40 909 -27
rect 943 -40 947 -27
rect 981 -40 985 -27
rect 1019 -40 1023 -27
rect 1057 -40 1061 -27
rect 1095 -40 1099 -27
rect 1133 -40 1137 -27
rect -17 -45 1161 -40
<< labels >>
rlabel metal1 -3 36 1 37 5 vdd
rlabel metal1 3 -42 7 -41 1 gnd
rlabel metal1 35 36 39 37 5 vdd
rlabel metal1 41 -42 45 -41 1 gnd
rlabel metal1 73 36 77 37 5 vdd
rlabel metal1 79 -42 83 -41 1 gnd
rlabel metal1 111 36 115 37 5 vdd
rlabel metal1 117 -42 121 -41 1 gnd
rlabel metal1 149 36 153 37 5 vdd
rlabel metal1 155 -42 159 -41 1 gnd
rlabel metal1 187 36 191 37 5 vdd
rlabel metal1 193 -42 197 -41 1 gnd
rlabel metal1 225 36 229 37 5 vdd
rlabel metal1 231 -42 235 -41 1 gnd
rlabel metal1 263 36 267 37 5 vdd
rlabel metal1 269 -42 273 -41 1 gnd
rlabel metal1 301 36 305 37 5 vdd
rlabel metal1 307 -42 311 -41 1 gnd
rlabel metal1 339 36 343 37 5 vdd
rlabel metal1 345 -42 349 -41 1 gnd
rlabel metal1 377 36 381 37 5 vdd
rlabel metal1 383 -42 387 -41 1 gnd
rlabel metal1 415 36 419 37 5 vdd
rlabel metal1 421 -42 425 -41 1 gnd
rlabel metal1 453 36 457 37 5 vdd
rlabel metal1 459 -42 463 -41 1 gnd
rlabel metal1 491 36 495 37 5 vdd
rlabel metal1 497 -42 501 -41 1 gnd
rlabel metal1 529 36 533 37 5 vdd
rlabel metal1 535 -42 539 -41 1 gnd
rlabel metal1 567 36 571 37 5 vdd
rlabel metal1 573 -42 577 -41 1 gnd
rlabel metal1 605 36 609 37 5 vdd
rlabel metal1 611 -42 615 -41 1 gnd
rlabel metal1 643 36 647 37 5 vdd
rlabel metal1 649 -42 653 -41 1 gnd
rlabel metal1 681 36 685 37 5 vdd
rlabel metal1 687 -42 691 -41 1 gnd
rlabel metal1 719 36 723 37 5 vdd
rlabel metal1 725 -42 729 -41 1 gnd
rlabel metal1 757 36 761 37 5 vdd
rlabel metal1 763 -42 767 -41 1 gnd
rlabel metal1 795 36 799 37 5 vdd
rlabel metal1 801 -42 805 -41 1 gnd
rlabel metal1 833 36 837 37 5 vdd
rlabel metal1 839 -42 843 -41 1 gnd
rlabel metal1 871 36 875 37 5 vdd
rlabel metal1 877 -42 881 -41 1 gnd
rlabel metal1 909 36 913 37 5 vdd
rlabel metal1 915 -42 919 -41 1 gnd
rlabel metal1 947 36 951 37 5 vdd
rlabel metal1 953 -42 957 -41 1 gnd
rlabel metal1 985 36 989 37 5 vdd
rlabel metal1 991 -42 995 -41 1 gnd
rlabel metal1 1023 36 1027 37 5 vdd
rlabel metal1 1029 -42 1033 -41 1 gnd
rlabel metal1 1061 36 1065 37 5 vdd
rlabel metal1 1067 -42 1071 -41 1 gnd
rlabel metal1 1099 36 1103 37 5 vdd
rlabel metal1 1105 -42 1109 -41 1 gnd
rlabel metal1 1137 36 1141 37 5 vdd
rlabel metal1 1143 -42 1147 -41 1 gnd
<< end >>
