.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.18u
.global gnd vdd

Vdd vdd gnd SUPPLY
vin a 0 pulse 0 1.8 0ns 100ps 100ps 9.9ns 20ns

.subckt inv y x vdd gnd
.param width_P={25*LAMBDA}
.param width_N={10*LAMBDA}
M1      y       x       gnd     gnd  CMOSN   W={width_N}   L={LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
M2      y       x       vdd     vdd  CMOSP   W={width_P}   L={LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
.ends inv

* inverter chain
x1 b a vdd gnd inv
x2 c b vdd gnd inv

Cload c gnd 100f   

.tran 0.1n 200n

.measure tran tpdr
+ TRIG v(a) VAL=SUPPLY/2 RISE=1
+ TARG v(c) VAL=SUPPLY/2 RISE=1

.measure tran tpdf
+ TRIG v(a) VAL=SUPPLY/2 FALL=1
+ TARG v(c) VAL=SUPPLY/2 FALL=1

.measure tran tpd param=(tpdr+tpdf)/2 goal=0

.control
set hcopypscolor = 1
set color0=white
set color1=black

run
plot v(a) v(c)
.endc
.end