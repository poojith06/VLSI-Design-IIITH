magic
tech scmos
timestamp 1764698600
<< nwell >>
rect -182 613 -120 621
rect -182 593 -69 613
rect -182 518 -120 526
rect -182 498 -69 518
rect 26 436 88 444
rect -181 422 -119 430
rect -181 402 -68 422
rect 26 416 139 436
rect 149 395 181 415
rect 193 395 225 415
rect 237 395 269 415
rect 281 395 313 415
rect 325 395 357 415
rect -177 328 -115 336
rect -177 308 -64 328
rect 5 301 25 337
rect 59 317 83 337
rect 3 277 25 301
rect 665 299 685 335
rect 739 326 801 334
rect 739 306 852 326
rect 663 275 685 299
rect -176 229 -114 237
rect 4 233 24 269
rect 54 253 78 273
rect -176 209 -63 229
rect 2 209 24 233
rect 665 224 685 260
rect 4 166 24 202
rect 54 186 78 206
rect 200 176 226 202
rect 247 176 273 202
rect 281 176 307 202
rect 328 176 354 202
rect 362 176 388 202
rect 409 176 435 202
rect 443 176 469 202
rect 490 176 516 202
rect 524 176 550 202
rect 571 176 597 202
rect 663 200 685 224
rect 739 231 801 239
rect 739 211 852 231
rect -175 153 -113 161
rect -175 133 -62 153
rect 2 142 24 166
rect 665 139 685 175
rect 4 96 24 132
rect 54 116 78 136
rect 663 115 685 139
rect 740 135 802 143
rect 740 115 853 135
rect 2 72 24 96
rect -180 49 -118 57
rect -180 29 -67 49
rect 4 24 24 60
rect 54 44 78 64
rect 674 52 694 88
rect 672 28 694 52
rect 744 41 806 49
rect 2 0 24 24
rect 744 21 857 41
rect -186 -65 -124 -57
rect -186 -85 -73 -65
rect 674 -84 694 -48
rect 745 -58 807 -50
rect 745 -78 858 -58
rect 672 -108 694 -84
rect 265 -142 297 -113
rect 319 -142 351 -113
rect 367 -142 399 -113
rect 415 -142 447 -113
rect 474 -142 506 -113
rect 747 -163 809 -155
rect 747 -183 860 -163
rect -189 -198 -127 -190
rect -189 -218 -76 -198
rect -190 -310 -128 -302
rect -190 -330 -77 -310
<< ntransistor >>
rect -171 581 -169 585
rect -141 579 -139 587
rect -133 579 -131 587
rect -106 576 -104 584
rect -98 576 -96 584
rect -82 581 -80 585
rect -171 486 -169 490
rect -141 484 -139 492
rect -133 484 -131 492
rect -106 481 -104 489
rect -98 481 -96 489
rect -82 486 -80 490
rect -170 390 -168 394
rect -140 388 -138 396
rect -132 388 -130 396
rect 37 404 39 408
rect 67 402 69 410
rect 75 402 77 410
rect -105 385 -103 393
rect -97 385 -95 393
rect -81 390 -79 394
rect 102 399 104 407
rect 110 399 112 407
rect 126 404 128 408
rect 160 375 162 383
rect 168 375 170 383
rect 204 375 206 383
rect 212 375 214 383
rect 248 375 250 383
rect 256 375 258 383
rect 292 375 294 383
rect 300 375 302 383
rect 336 375 338 383
rect 344 375 346 383
rect 31 324 35 326
rect -166 296 -164 300
rect -136 294 -134 302
rect -128 294 -126 302
rect 31 306 35 308
rect 691 322 695 324
rect 70 302 72 306
rect 691 304 695 306
rect -101 291 -99 299
rect -93 291 -91 299
rect -77 296 -75 300
rect 750 294 752 298
rect 35 288 39 290
rect 780 292 782 300
rect 788 292 790 300
rect 695 286 699 288
rect 815 289 817 297
rect 823 289 825 297
rect 839 294 841 298
rect 30 256 34 258
rect 691 247 695 249
rect 30 238 34 240
rect 65 238 67 242
rect 691 229 695 231
rect 34 220 38 222
rect -165 197 -163 201
rect -135 195 -133 203
rect -127 195 -125 203
rect 695 211 699 213
rect -100 192 -98 200
rect -92 192 -90 200
rect -76 197 -74 201
rect 750 199 752 203
rect 30 189 34 191
rect 780 197 782 205
rect 788 197 790 205
rect 815 194 817 202
rect 823 194 825 202
rect 839 199 841 203
rect 30 171 34 173
rect 65 171 67 175
rect 212 162 214 166
rect 34 153 38 155
rect 259 161 261 165
rect 293 162 295 166
rect 340 161 342 165
rect 374 162 376 166
rect 421 161 423 165
rect 455 162 457 166
rect 502 161 504 165
rect 536 162 538 166
rect 583 161 585 165
rect 691 162 695 164
rect 691 144 695 146
rect -164 121 -162 125
rect -134 119 -132 127
rect -126 119 -124 127
rect -99 116 -97 124
rect -91 116 -89 124
rect -75 121 -73 125
rect 695 126 699 128
rect 30 119 34 121
rect 30 101 34 103
rect 65 101 67 105
rect 751 103 753 107
rect 781 101 783 109
rect 789 101 791 109
rect 816 98 818 106
rect 824 98 826 106
rect 840 103 842 107
rect 34 83 38 85
rect 700 75 704 77
rect 700 57 704 59
rect 30 47 34 49
rect -169 17 -167 21
rect -139 15 -137 23
rect -131 15 -129 23
rect 704 39 708 41
rect 30 29 34 31
rect 65 29 67 33
rect -104 12 -102 20
rect -96 12 -94 20
rect -80 17 -78 21
rect 34 11 38 13
rect 755 9 757 13
rect 785 7 787 15
rect 793 7 795 15
rect 820 4 822 12
rect 828 4 830 12
rect 844 9 846 13
rect 700 -61 704 -59
rect 700 -79 704 -77
rect -175 -97 -173 -93
rect -145 -99 -143 -91
rect -137 -99 -135 -91
rect 756 -90 758 -86
rect -110 -102 -108 -94
rect -102 -102 -100 -94
rect -86 -97 -84 -93
rect 786 -92 788 -84
rect 794 -92 796 -84
rect 704 -97 708 -95
rect 276 -104 278 -100
rect 284 -104 286 -100
rect 330 -104 332 -100
rect 338 -104 340 -100
rect 378 -104 380 -100
rect 386 -104 388 -100
rect 426 -104 428 -100
rect 434 -104 436 -100
rect 485 -104 487 -100
rect 493 -104 495 -100
rect 821 -95 823 -87
rect 829 -95 831 -87
rect 845 -90 847 -86
rect 758 -195 760 -191
rect 788 -197 790 -189
rect 796 -197 798 -189
rect 823 -200 825 -192
rect 831 -200 833 -192
rect 847 -195 849 -191
rect -178 -230 -176 -226
rect -148 -232 -146 -224
rect -140 -232 -138 -224
rect -113 -235 -111 -227
rect -105 -235 -103 -227
rect -89 -230 -87 -226
rect -179 -342 -177 -338
rect -149 -344 -147 -336
rect -141 -344 -139 -336
rect -114 -347 -112 -339
rect -106 -347 -104 -339
rect -90 -342 -88 -338
<< ptransistor >>
rect -171 599 -169 615
rect -163 599 -161 615
rect -141 599 -139 615
rect -133 599 -131 615
rect -116 599 -114 607
rect -98 599 -96 607
rect -82 599 -80 607
rect -171 504 -169 520
rect -163 504 -161 520
rect -141 504 -139 520
rect -133 504 -131 520
rect -116 504 -114 512
rect -98 504 -96 512
rect -82 504 -80 512
rect -170 408 -168 424
rect -162 408 -160 424
rect -140 408 -138 424
rect -132 408 -130 424
rect 37 422 39 438
rect 45 422 47 438
rect 67 422 69 438
rect 75 422 77 438
rect 92 422 94 430
rect 110 422 112 430
rect 126 422 128 430
rect -115 408 -113 416
rect -97 408 -95 416
rect -81 408 -79 416
rect 160 401 162 409
rect 168 401 170 409
rect 204 401 206 409
rect 212 401 214 409
rect 248 401 250 409
rect 256 401 258 409
rect 292 401 294 409
rect 300 401 302 409
rect 336 401 338 409
rect 344 401 346 409
rect -166 314 -164 330
rect -158 314 -156 330
rect -136 314 -134 330
rect -128 314 -126 330
rect 11 324 19 326
rect -111 314 -109 322
rect -93 314 -91 322
rect -77 314 -75 322
rect 70 323 72 331
rect 11 306 19 308
rect 671 322 679 324
rect 750 312 752 328
rect 758 312 760 328
rect 780 312 782 328
rect 788 312 790 328
rect 805 312 807 320
rect 823 312 825 320
rect 839 312 841 320
rect 671 304 679 306
rect 11 288 19 290
rect 671 286 679 288
rect 65 259 67 267
rect 10 256 18 258
rect 671 247 679 249
rect 10 238 18 240
rect -165 215 -163 231
rect -157 215 -155 231
rect -135 215 -133 231
rect -127 215 -125 231
rect 671 229 679 231
rect -110 215 -108 223
rect -92 215 -90 223
rect -76 215 -74 223
rect 10 220 18 222
rect 750 217 752 233
rect 758 217 760 233
rect 780 217 782 233
rect 788 217 790 233
rect 805 217 807 225
rect 823 217 825 225
rect 839 217 841 225
rect 671 211 679 213
rect 65 192 67 200
rect 10 189 18 191
rect 212 183 214 191
rect 259 183 261 191
rect 293 183 295 191
rect 340 183 342 191
rect 374 183 376 191
rect 421 183 423 191
rect 455 183 457 191
rect 502 183 504 191
rect 536 183 538 191
rect 583 183 585 191
rect 10 171 18 173
rect -164 139 -162 155
rect -156 139 -154 155
rect -134 139 -132 155
rect -126 139 -124 155
rect 10 153 18 155
rect 671 162 679 164
rect -109 139 -107 147
rect -91 139 -89 147
rect -75 139 -73 147
rect 671 144 679 146
rect 65 122 67 130
rect 671 126 679 128
rect 10 119 18 121
rect 751 121 753 137
rect 759 121 761 137
rect 781 121 783 137
rect 789 121 791 137
rect 806 121 808 129
rect 824 121 826 129
rect 840 121 842 129
rect 10 101 18 103
rect 10 83 18 85
rect 680 75 688 77
rect -169 35 -167 51
rect -161 35 -159 51
rect -139 35 -137 51
rect -131 35 -129 51
rect 65 50 67 58
rect 680 57 688 59
rect 10 47 18 49
rect -114 35 -112 43
rect -96 35 -94 43
rect -80 35 -78 43
rect 680 39 688 41
rect 10 29 18 31
rect 755 27 757 43
rect 763 27 765 43
rect 785 27 787 43
rect 793 27 795 43
rect 810 27 812 35
rect 828 27 830 35
rect 844 27 846 35
rect 10 11 18 13
rect -175 -79 -173 -63
rect -167 -79 -165 -63
rect -145 -79 -143 -63
rect -137 -79 -135 -63
rect 680 -61 688 -59
rect -120 -79 -118 -71
rect -102 -79 -100 -71
rect -86 -79 -84 -71
rect 756 -72 758 -56
rect 764 -72 766 -56
rect 786 -72 788 -56
rect 794 -72 796 -56
rect 811 -72 813 -64
rect 829 -72 831 -64
rect 845 -72 847 -64
rect 680 -79 688 -77
rect 680 -97 688 -95
rect 276 -136 278 -120
rect 284 -136 286 -120
rect 330 -136 332 -120
rect 338 -136 340 -120
rect 378 -136 380 -120
rect 386 -136 388 -120
rect 426 -136 428 -120
rect 434 -136 436 -120
rect 485 -136 487 -120
rect 493 -136 495 -120
rect 758 -177 760 -161
rect 766 -177 768 -161
rect 788 -177 790 -161
rect 796 -177 798 -161
rect 813 -177 815 -169
rect 831 -177 833 -169
rect 847 -177 849 -169
rect -178 -212 -176 -196
rect -170 -212 -168 -196
rect -148 -212 -146 -196
rect -140 -212 -138 -196
rect -123 -212 -121 -204
rect -105 -212 -103 -204
rect -89 -212 -87 -204
rect -179 -324 -177 -308
rect -171 -324 -169 -308
rect -149 -324 -147 -308
rect -141 -324 -139 -308
rect -124 -324 -122 -316
rect -106 -324 -104 -316
rect -90 -324 -88 -316
<< ndiffusion >>
rect -172 581 -171 585
rect -169 581 -168 585
rect -142 579 -141 587
rect -139 579 -138 587
rect -134 579 -133 587
rect -131 579 -130 587
rect -107 576 -106 584
rect -104 576 -103 584
rect -99 576 -98 584
rect -96 576 -95 584
rect -83 581 -82 585
rect -80 581 -79 585
rect -172 486 -171 490
rect -169 486 -168 490
rect -142 484 -141 492
rect -139 484 -138 492
rect -134 484 -133 492
rect -131 484 -130 492
rect -107 481 -106 489
rect -104 481 -103 489
rect -99 481 -98 489
rect -96 481 -95 489
rect -83 486 -82 490
rect -80 486 -79 490
rect -171 390 -170 394
rect -168 390 -167 394
rect -141 388 -140 396
rect -138 388 -137 396
rect -133 388 -132 396
rect -130 388 -129 396
rect 36 404 37 408
rect 39 404 40 408
rect 66 402 67 410
rect 69 402 70 410
rect 74 402 75 410
rect 77 402 78 410
rect -106 385 -105 393
rect -103 385 -102 393
rect -98 385 -97 393
rect -95 385 -94 393
rect -82 390 -81 394
rect -79 390 -78 394
rect 101 399 102 407
rect 104 399 105 407
rect 109 399 110 407
rect 112 399 113 407
rect 125 404 126 408
rect 128 404 129 408
rect 159 375 160 383
rect 162 375 163 383
rect 167 375 168 383
rect 170 375 171 383
rect 203 375 204 383
rect 206 375 207 383
rect 211 375 212 383
rect 214 375 215 383
rect 247 375 248 383
rect 250 375 251 383
rect 255 375 256 383
rect 258 375 259 383
rect 291 375 292 383
rect 294 375 295 383
rect 299 375 300 383
rect 302 375 303 383
rect 335 375 336 383
rect 338 375 339 383
rect 343 375 344 383
rect 346 375 347 383
rect 31 326 35 327
rect 31 323 35 324
rect 691 324 695 325
rect -167 296 -166 300
rect -164 296 -163 300
rect -137 294 -136 302
rect -134 294 -133 302
rect -129 294 -128 302
rect -126 294 -125 302
rect 31 308 35 309
rect 691 321 695 322
rect 691 306 695 307
rect 31 305 35 306
rect 69 302 70 306
rect 72 302 73 306
rect -102 291 -101 299
rect -99 291 -98 299
rect -94 291 -93 299
rect -91 291 -90 299
rect -78 296 -77 300
rect -75 296 -74 300
rect 691 303 695 304
rect 749 294 750 298
rect 752 294 753 298
rect 35 290 39 291
rect 779 292 780 300
rect 782 292 783 300
rect 787 292 788 300
rect 790 292 791 300
rect 695 288 699 289
rect 35 287 39 288
rect 695 285 699 286
rect 814 289 815 297
rect 817 289 818 297
rect 822 289 823 297
rect 825 289 826 297
rect 838 294 839 298
rect 841 294 842 298
rect 30 258 34 259
rect 30 255 34 256
rect 691 249 695 250
rect 691 246 695 247
rect 30 240 34 241
rect 64 238 65 242
rect 67 238 68 242
rect 30 237 34 238
rect 691 231 695 232
rect 691 228 695 229
rect 34 222 38 223
rect 34 219 38 220
rect -166 197 -165 201
rect -163 197 -162 201
rect -136 195 -135 203
rect -133 195 -132 203
rect -128 195 -127 203
rect -125 195 -124 203
rect 695 213 699 214
rect 695 210 699 211
rect -101 192 -100 200
rect -98 192 -97 200
rect -93 192 -92 200
rect -90 192 -89 200
rect -77 197 -76 201
rect -74 197 -73 201
rect 749 199 750 203
rect 752 199 753 203
rect 30 191 34 192
rect 30 188 34 189
rect 779 197 780 205
rect 782 197 783 205
rect 787 197 788 205
rect 790 197 791 205
rect 814 194 815 202
rect 817 194 818 202
rect 822 194 823 202
rect 825 194 826 202
rect 838 199 839 203
rect 841 199 842 203
rect 30 173 34 174
rect 64 171 65 175
rect 67 171 68 175
rect 30 170 34 171
rect 211 162 212 166
rect 214 162 215 166
rect 34 155 38 156
rect 34 152 38 153
rect 258 161 259 165
rect 261 161 262 165
rect 292 162 293 166
rect 295 162 296 166
rect 339 161 340 165
rect 342 161 343 165
rect 373 162 374 166
rect 376 162 377 166
rect 420 161 421 165
rect 423 161 424 165
rect 454 162 455 166
rect 457 162 458 166
rect 501 161 502 165
rect 504 161 505 165
rect 535 162 536 166
rect 538 162 539 166
rect 582 161 583 165
rect 585 161 586 165
rect 691 164 695 165
rect 691 161 695 162
rect 691 146 695 147
rect 691 143 695 144
rect -165 121 -164 125
rect -162 121 -161 125
rect -135 119 -134 127
rect -132 119 -131 127
rect -127 119 -126 127
rect -124 119 -123 127
rect -100 116 -99 124
rect -97 116 -96 124
rect -92 116 -91 124
rect -89 116 -88 124
rect -76 121 -75 125
rect -73 121 -72 125
rect 695 128 699 129
rect 30 121 34 122
rect 30 118 34 119
rect 695 125 699 126
rect 30 103 34 104
rect 64 101 65 105
rect 67 101 68 105
rect 750 103 751 107
rect 753 103 754 107
rect 30 100 34 101
rect 780 101 781 109
rect 783 101 784 109
rect 788 101 789 109
rect 791 101 792 109
rect 815 98 816 106
rect 818 98 819 106
rect 823 98 824 106
rect 826 98 827 106
rect 839 103 840 107
rect 842 103 843 107
rect 34 85 38 86
rect 34 82 38 83
rect 700 77 704 78
rect 700 74 704 75
rect 700 59 704 60
rect 700 56 704 57
rect 30 49 34 50
rect 30 46 34 47
rect -170 17 -169 21
rect -167 17 -166 21
rect -140 15 -139 23
rect -137 15 -136 23
rect -132 15 -131 23
rect -129 15 -128 23
rect 704 41 708 42
rect 704 38 708 39
rect 30 31 34 32
rect 64 29 65 33
rect 67 29 68 33
rect 30 28 34 29
rect -105 12 -104 20
rect -102 12 -101 20
rect -97 12 -96 20
rect -94 12 -93 20
rect -81 17 -80 21
rect -78 17 -77 21
rect 34 13 38 14
rect 34 10 38 11
rect 754 9 755 13
rect 757 9 758 13
rect 784 7 785 15
rect 787 7 788 15
rect 792 7 793 15
rect 795 7 796 15
rect 819 4 820 12
rect 822 4 823 12
rect 827 4 828 12
rect 830 4 831 12
rect 843 9 844 13
rect 846 9 847 13
rect 700 -59 704 -58
rect 700 -62 704 -61
rect 700 -77 704 -76
rect -176 -97 -175 -93
rect -173 -97 -172 -93
rect -146 -99 -145 -91
rect -143 -99 -142 -91
rect -138 -99 -137 -91
rect -135 -99 -134 -91
rect 700 -80 704 -79
rect 755 -90 756 -86
rect 758 -90 759 -86
rect -111 -102 -110 -94
rect -108 -102 -107 -94
rect -103 -102 -102 -94
rect -100 -102 -99 -94
rect -87 -97 -86 -93
rect -84 -97 -83 -93
rect 785 -92 786 -84
rect 788 -92 789 -84
rect 793 -92 794 -84
rect 796 -92 797 -84
rect 704 -95 708 -94
rect 275 -104 276 -100
rect 278 -104 279 -100
rect 283 -104 284 -100
rect 286 -104 287 -100
rect 329 -104 330 -100
rect 332 -104 333 -100
rect 337 -104 338 -100
rect 340 -104 341 -100
rect 377 -104 378 -100
rect 380 -104 381 -100
rect 385 -104 386 -100
rect 388 -104 389 -100
rect 425 -104 426 -100
rect 428 -104 429 -100
rect 433 -104 434 -100
rect 436 -104 437 -100
rect 484 -104 485 -100
rect 487 -104 488 -100
rect 492 -104 493 -100
rect 495 -104 496 -100
rect 704 -98 708 -97
rect 820 -95 821 -87
rect 823 -95 824 -87
rect 828 -95 829 -87
rect 831 -95 832 -87
rect 844 -90 845 -86
rect 847 -90 848 -86
rect 757 -195 758 -191
rect 760 -195 761 -191
rect 787 -197 788 -189
rect 790 -197 791 -189
rect 795 -197 796 -189
rect 798 -197 799 -189
rect 822 -200 823 -192
rect 825 -200 826 -192
rect 830 -200 831 -192
rect 833 -200 834 -192
rect 846 -195 847 -191
rect 849 -195 850 -191
rect -179 -230 -178 -226
rect -176 -230 -175 -226
rect -149 -232 -148 -224
rect -146 -232 -145 -224
rect -141 -232 -140 -224
rect -138 -232 -137 -224
rect -114 -235 -113 -227
rect -111 -235 -110 -227
rect -106 -235 -105 -227
rect -103 -235 -102 -227
rect -90 -230 -89 -226
rect -87 -230 -86 -226
rect -180 -342 -179 -338
rect -177 -342 -176 -338
rect -150 -344 -149 -336
rect -147 -344 -146 -336
rect -142 -344 -141 -336
rect -139 -344 -138 -336
rect -115 -347 -114 -339
rect -112 -347 -111 -339
rect -107 -347 -106 -339
rect -104 -347 -103 -339
rect -91 -342 -90 -338
rect -88 -342 -87 -338
<< pdiffusion >>
rect -172 599 -171 615
rect -169 599 -168 615
rect -164 599 -163 615
rect -161 599 -160 615
rect -142 599 -141 615
rect -139 599 -138 615
rect -134 599 -133 615
rect -131 599 -130 615
rect -117 599 -116 607
rect -114 599 -113 607
rect -99 599 -98 607
rect -96 599 -95 607
rect -83 599 -82 607
rect -80 599 -79 607
rect -172 504 -171 520
rect -169 504 -168 520
rect -164 504 -163 520
rect -161 504 -160 520
rect -142 504 -141 520
rect -139 504 -138 520
rect -134 504 -133 520
rect -131 504 -130 520
rect -117 504 -116 512
rect -114 504 -113 512
rect -99 504 -98 512
rect -96 504 -95 512
rect -83 504 -82 512
rect -80 504 -79 512
rect -171 408 -170 424
rect -168 408 -167 424
rect -163 408 -162 424
rect -160 408 -159 424
rect -141 408 -140 424
rect -138 408 -137 424
rect -133 408 -132 424
rect -130 408 -129 424
rect 36 422 37 438
rect 39 422 40 438
rect 44 422 45 438
rect 47 422 48 438
rect 66 422 67 438
rect 69 422 70 438
rect 74 422 75 438
rect 77 422 78 438
rect 91 422 92 430
rect 94 422 95 430
rect 109 422 110 430
rect 112 422 113 430
rect 125 422 126 430
rect 128 422 129 430
rect -116 408 -115 416
rect -113 408 -112 416
rect -98 408 -97 416
rect -95 408 -94 416
rect -82 408 -81 416
rect -79 408 -78 416
rect 159 401 160 409
rect 162 401 163 409
rect 167 401 168 409
rect 170 401 171 409
rect 203 401 204 409
rect 206 401 207 409
rect 211 401 212 409
rect 214 401 215 409
rect 247 401 248 409
rect 250 401 251 409
rect 255 401 256 409
rect 258 401 259 409
rect 291 401 292 409
rect 294 401 295 409
rect 299 401 300 409
rect 302 401 303 409
rect 335 401 336 409
rect 338 401 339 409
rect 343 401 344 409
rect 346 401 347 409
rect -167 314 -166 330
rect -164 314 -163 330
rect -159 314 -158 330
rect -156 314 -155 330
rect -137 314 -136 330
rect -134 314 -133 330
rect -129 314 -128 330
rect -126 314 -125 330
rect 11 326 19 327
rect -112 314 -111 322
rect -109 314 -108 322
rect -94 314 -93 322
rect -91 314 -90 322
rect -78 314 -77 322
rect -75 314 -74 322
rect 11 323 19 324
rect 69 323 70 331
rect 72 323 73 331
rect 671 324 679 325
rect 11 308 19 309
rect 671 321 679 322
rect 749 312 750 328
rect 752 312 753 328
rect 757 312 758 328
rect 760 312 761 328
rect 779 312 780 328
rect 782 312 783 328
rect 787 312 788 328
rect 790 312 791 328
rect 804 312 805 320
rect 807 312 808 320
rect 822 312 823 320
rect 825 312 826 320
rect 838 312 839 320
rect 841 312 842 320
rect 671 306 679 307
rect 11 305 19 306
rect 671 303 679 304
rect 11 290 19 291
rect 671 288 679 289
rect 11 287 19 288
rect 671 285 679 286
rect 10 258 18 259
rect 64 259 65 267
rect 67 259 68 267
rect 10 255 18 256
rect 10 240 18 241
rect 671 249 679 250
rect 671 246 679 247
rect 10 237 18 238
rect -166 215 -165 231
rect -163 215 -162 231
rect -158 215 -157 231
rect -155 215 -154 231
rect -136 215 -135 231
rect -133 215 -132 231
rect -128 215 -127 231
rect -125 215 -124 231
rect 671 231 679 232
rect 671 228 679 229
rect -111 215 -110 223
rect -108 215 -107 223
rect -93 215 -92 223
rect -90 215 -89 223
rect -77 215 -76 223
rect -74 215 -73 223
rect 10 222 18 223
rect 10 219 18 220
rect 671 213 679 214
rect 749 217 750 233
rect 752 217 753 233
rect 757 217 758 233
rect 760 217 761 233
rect 779 217 780 233
rect 782 217 783 233
rect 787 217 788 233
rect 790 217 791 233
rect 804 217 805 225
rect 807 217 808 225
rect 822 217 823 225
rect 825 217 826 225
rect 838 217 839 225
rect 841 217 842 225
rect 671 210 679 211
rect 10 191 18 192
rect 64 192 65 200
rect 67 192 68 200
rect 10 188 18 189
rect 10 173 18 174
rect 211 183 212 191
rect 214 183 215 191
rect 258 183 259 191
rect 261 183 262 191
rect 292 183 293 191
rect 295 183 296 191
rect 339 183 340 191
rect 342 183 343 191
rect 373 183 374 191
rect 376 183 377 191
rect 420 183 421 191
rect 423 183 424 191
rect 454 183 455 191
rect 457 183 458 191
rect 501 183 502 191
rect 504 183 505 191
rect 535 183 536 191
rect 538 183 539 191
rect 582 183 583 191
rect 585 183 586 191
rect 10 170 18 171
rect -165 139 -164 155
rect -162 139 -161 155
rect -157 139 -156 155
rect -154 139 -153 155
rect -135 139 -134 155
rect -132 139 -131 155
rect -127 139 -126 155
rect -124 139 -123 155
rect 10 155 18 156
rect 10 152 18 153
rect 671 164 679 165
rect 671 161 679 162
rect -110 139 -109 147
rect -107 139 -106 147
rect -92 139 -91 147
rect -89 139 -88 147
rect -76 139 -75 147
rect -73 139 -72 147
rect 671 146 679 147
rect 671 143 679 144
rect 10 121 18 122
rect 64 122 65 130
rect 67 122 68 130
rect 671 128 679 129
rect 671 125 679 126
rect 10 118 18 119
rect 10 103 18 104
rect 750 121 751 137
rect 753 121 754 137
rect 758 121 759 137
rect 761 121 762 137
rect 780 121 781 137
rect 783 121 784 137
rect 788 121 789 137
rect 791 121 792 137
rect 805 121 806 129
rect 808 121 809 129
rect 823 121 824 129
rect 826 121 827 129
rect 839 121 840 129
rect 842 121 843 129
rect 10 100 18 101
rect 10 85 18 86
rect 10 82 18 83
rect 680 77 688 78
rect 680 74 688 75
rect 680 59 688 60
rect -170 35 -169 51
rect -167 35 -166 51
rect -162 35 -161 51
rect -159 35 -158 51
rect -140 35 -139 51
rect -137 35 -136 51
rect -132 35 -131 51
rect -129 35 -128 51
rect 10 49 18 50
rect 64 50 65 58
rect 67 50 68 58
rect 680 56 688 57
rect 10 46 18 47
rect -115 35 -114 43
rect -112 35 -111 43
rect -97 35 -96 43
rect -94 35 -93 43
rect -81 35 -80 43
rect -78 35 -77 43
rect 10 31 18 32
rect 680 41 688 42
rect 680 38 688 39
rect 10 28 18 29
rect 754 27 755 43
rect 757 27 758 43
rect 762 27 763 43
rect 765 27 766 43
rect 784 27 785 43
rect 787 27 788 43
rect 792 27 793 43
rect 795 27 796 43
rect 809 27 810 35
rect 812 27 813 35
rect 827 27 828 35
rect 830 27 831 35
rect 843 27 844 35
rect 846 27 847 35
rect 10 13 18 14
rect 10 10 18 11
rect -176 -79 -175 -63
rect -173 -79 -172 -63
rect -168 -79 -167 -63
rect -165 -79 -164 -63
rect -146 -79 -145 -63
rect -143 -79 -142 -63
rect -138 -79 -137 -63
rect -135 -79 -134 -63
rect 680 -59 688 -58
rect 680 -62 688 -61
rect -121 -79 -120 -71
rect -118 -79 -117 -71
rect -103 -79 -102 -71
rect -100 -79 -99 -71
rect -87 -79 -86 -71
rect -84 -79 -83 -71
rect 755 -72 756 -56
rect 758 -72 759 -56
rect 763 -72 764 -56
rect 766 -72 767 -56
rect 785 -72 786 -56
rect 788 -72 789 -56
rect 793 -72 794 -56
rect 796 -72 797 -56
rect 810 -72 811 -64
rect 813 -72 814 -64
rect 828 -72 829 -64
rect 831 -72 832 -64
rect 844 -72 845 -64
rect 847 -72 848 -64
rect 680 -77 688 -76
rect 680 -80 688 -79
rect 680 -95 688 -94
rect 680 -98 688 -97
rect 275 -136 276 -120
rect 278 -136 279 -120
rect 283 -136 284 -120
rect 286 -136 287 -120
rect 329 -136 330 -120
rect 332 -136 333 -120
rect 337 -136 338 -120
rect 340 -136 341 -120
rect 377 -136 378 -120
rect 380 -136 381 -120
rect 385 -136 386 -120
rect 388 -136 389 -120
rect 425 -136 426 -120
rect 428 -136 429 -120
rect 433 -136 434 -120
rect 436 -136 437 -120
rect 484 -136 485 -120
rect 487 -136 488 -120
rect 492 -136 493 -120
rect 495 -136 496 -120
rect 757 -177 758 -161
rect 760 -177 761 -161
rect 765 -177 766 -161
rect 768 -177 769 -161
rect 787 -177 788 -161
rect 790 -177 791 -161
rect 795 -177 796 -161
rect 798 -177 799 -161
rect 812 -177 813 -169
rect 815 -177 816 -169
rect 830 -177 831 -169
rect 833 -177 834 -169
rect 846 -177 847 -169
rect 849 -177 850 -169
rect -179 -212 -178 -196
rect -176 -212 -175 -196
rect -171 -212 -170 -196
rect -168 -212 -167 -196
rect -149 -212 -148 -196
rect -146 -212 -145 -196
rect -141 -212 -140 -196
rect -138 -212 -137 -196
rect -124 -212 -123 -204
rect -121 -212 -120 -204
rect -106 -212 -105 -204
rect -103 -212 -102 -204
rect -90 -212 -89 -204
rect -87 -212 -86 -204
rect -180 -324 -179 -308
rect -177 -324 -176 -308
rect -172 -324 -171 -308
rect -169 -324 -168 -308
rect -150 -324 -149 -308
rect -147 -324 -146 -308
rect -142 -324 -141 -308
rect -139 -324 -138 -308
rect -125 -324 -124 -316
rect -122 -324 -121 -316
rect -107 -324 -106 -316
rect -104 -324 -103 -316
rect -91 -324 -90 -316
rect -88 -324 -87 -316
<< ndcontact >>
rect -176 581 -172 585
rect -168 581 -164 585
rect -146 579 -142 587
rect -138 579 -134 587
rect -130 579 -126 587
rect -111 576 -107 584
rect -103 576 -99 584
rect -95 576 -91 584
rect -87 581 -83 585
rect -79 581 -75 585
rect -176 486 -172 490
rect -168 486 -164 490
rect -146 484 -142 492
rect -138 484 -134 492
rect -130 484 -126 492
rect -111 481 -107 489
rect -103 481 -99 489
rect -95 481 -91 489
rect -87 486 -83 490
rect -79 486 -75 490
rect -175 390 -171 394
rect -167 390 -163 394
rect -145 388 -141 396
rect -137 388 -133 396
rect -129 388 -125 396
rect 32 404 36 408
rect 40 404 44 408
rect 62 402 66 410
rect 70 402 74 410
rect 78 402 82 410
rect -110 385 -106 393
rect -102 385 -98 393
rect -94 385 -90 393
rect -86 390 -82 394
rect -78 390 -74 394
rect 97 399 101 407
rect 105 399 109 407
rect 113 399 117 407
rect 121 404 125 408
rect 129 404 133 408
rect 155 375 159 383
rect 163 375 167 383
rect 171 375 175 383
rect 199 375 203 383
rect 207 375 211 383
rect 215 375 219 383
rect 243 375 247 383
rect 251 375 255 383
rect 259 375 263 383
rect 287 375 291 383
rect 295 375 299 383
rect 303 375 307 383
rect 331 375 335 383
rect 339 375 343 383
rect 347 375 351 383
rect 31 327 35 331
rect 31 319 35 323
rect 691 325 695 329
rect -171 296 -167 300
rect -163 296 -159 300
rect -141 294 -137 302
rect -133 294 -129 302
rect -125 294 -121 302
rect 31 309 35 313
rect 691 317 695 321
rect 691 307 695 311
rect 31 301 35 305
rect 65 302 69 306
rect 73 302 77 306
rect -106 291 -102 299
rect -98 291 -94 299
rect -90 291 -86 299
rect -82 296 -78 300
rect -74 296 -70 300
rect 691 299 695 303
rect 35 291 39 295
rect 745 294 749 298
rect 753 294 757 298
rect 695 289 699 293
rect 775 292 779 300
rect 783 292 787 300
rect 791 292 795 300
rect 35 283 39 287
rect 695 281 699 285
rect 810 289 814 297
rect 818 289 822 297
rect 826 289 830 297
rect 834 294 838 298
rect 842 294 846 298
rect 30 259 34 263
rect 30 251 34 255
rect 30 241 34 245
rect 691 250 695 254
rect 691 242 695 246
rect 60 238 64 242
rect 68 238 72 242
rect 30 233 34 237
rect 691 232 695 236
rect 34 223 38 227
rect 691 224 695 228
rect 34 215 38 219
rect -170 197 -166 201
rect -162 197 -158 201
rect -140 195 -136 203
rect -132 195 -128 203
rect -124 195 -120 203
rect 695 214 699 218
rect 695 206 699 210
rect -105 192 -101 200
rect -97 192 -93 200
rect -89 192 -85 200
rect -81 197 -77 201
rect -73 197 -69 201
rect 30 192 34 196
rect 745 199 749 203
rect 753 199 757 203
rect 30 184 34 188
rect 30 174 34 178
rect 775 197 779 205
rect 783 197 787 205
rect 791 197 795 205
rect 810 194 814 202
rect 818 194 822 202
rect 826 194 830 202
rect 834 199 838 203
rect 842 199 846 203
rect 60 171 64 175
rect 68 171 72 175
rect 30 166 34 170
rect 207 162 211 166
rect 215 162 219 166
rect 34 156 38 160
rect 254 161 258 165
rect 262 161 266 165
rect 288 162 292 166
rect 296 162 300 166
rect 335 161 339 165
rect 343 161 347 165
rect 369 162 373 166
rect 377 162 381 166
rect 416 161 420 165
rect 424 161 428 165
rect 450 162 454 166
rect 458 162 462 166
rect 497 161 501 165
rect 505 161 509 165
rect 531 162 535 166
rect 539 162 543 166
rect 578 161 582 165
rect 586 161 590 165
rect 691 165 695 169
rect 691 157 695 161
rect 34 148 38 152
rect 691 147 695 151
rect 691 139 695 143
rect -169 121 -165 125
rect -161 121 -157 125
rect -139 119 -135 127
rect -131 119 -127 127
rect -123 119 -119 127
rect -104 116 -100 124
rect -96 116 -92 124
rect -88 116 -84 124
rect -80 121 -76 125
rect -72 121 -68 125
rect 30 122 34 126
rect 695 129 699 133
rect 30 114 34 118
rect 30 104 34 108
rect 695 121 699 125
rect 60 101 64 105
rect 68 101 72 105
rect 746 103 750 107
rect 754 103 758 107
rect 30 96 34 100
rect 776 101 780 109
rect 784 101 788 109
rect 792 101 796 109
rect 811 98 815 106
rect 819 98 823 106
rect 827 98 831 106
rect 835 103 839 107
rect 843 103 847 107
rect 34 86 38 90
rect 34 78 38 82
rect 700 78 704 82
rect 700 70 704 74
rect 700 60 704 64
rect 30 50 34 54
rect 700 52 704 56
rect 30 42 34 46
rect -174 17 -170 21
rect -166 17 -162 21
rect -144 15 -140 23
rect -136 15 -132 23
rect -128 15 -124 23
rect 30 32 34 36
rect 704 42 708 46
rect 704 34 708 38
rect 60 29 64 33
rect 68 29 72 33
rect 30 24 34 28
rect -109 12 -105 20
rect -101 12 -97 20
rect -93 12 -89 20
rect -85 17 -81 21
rect -77 17 -73 21
rect 34 14 38 18
rect 34 6 38 10
rect 750 9 754 13
rect 758 9 762 13
rect 780 7 784 15
rect 788 7 792 15
rect 796 7 800 15
rect 815 4 819 12
rect 823 4 827 12
rect 831 4 835 12
rect 839 9 843 13
rect 847 9 851 13
rect 700 -58 704 -54
rect 700 -66 704 -62
rect 700 -76 704 -72
rect -180 -97 -176 -93
rect -172 -97 -168 -93
rect -150 -99 -146 -91
rect -142 -99 -138 -91
rect -134 -99 -130 -91
rect 700 -84 704 -80
rect 751 -90 755 -86
rect 759 -90 763 -86
rect -115 -102 -111 -94
rect -107 -102 -103 -94
rect -99 -102 -95 -94
rect -91 -97 -87 -93
rect -83 -97 -79 -93
rect 704 -94 708 -90
rect 781 -92 785 -84
rect 789 -92 793 -84
rect 797 -92 801 -84
rect 271 -104 275 -100
rect 279 -104 283 -100
rect 287 -104 291 -100
rect 325 -104 329 -100
rect 333 -104 337 -100
rect 341 -104 345 -100
rect 373 -104 377 -100
rect 381 -104 385 -100
rect 389 -104 393 -100
rect 421 -104 425 -100
rect 429 -104 433 -100
rect 437 -104 441 -100
rect 480 -104 484 -100
rect 488 -104 492 -100
rect 496 -104 500 -100
rect 704 -102 708 -98
rect 816 -95 820 -87
rect 824 -95 828 -87
rect 832 -95 836 -87
rect 840 -90 844 -86
rect 848 -90 852 -86
rect 753 -195 757 -191
rect 761 -195 765 -191
rect 783 -197 787 -189
rect 791 -197 795 -189
rect 799 -197 803 -189
rect 818 -200 822 -192
rect 826 -200 830 -192
rect 834 -200 838 -192
rect 842 -195 846 -191
rect 850 -195 854 -191
rect -183 -230 -179 -226
rect -175 -230 -171 -226
rect -153 -232 -149 -224
rect -145 -232 -141 -224
rect -137 -232 -133 -224
rect -118 -235 -114 -227
rect -110 -235 -106 -227
rect -102 -235 -98 -227
rect -94 -230 -90 -226
rect -86 -230 -82 -226
rect -184 -342 -180 -338
rect -176 -342 -172 -338
rect -154 -344 -150 -336
rect -146 -344 -142 -336
rect -138 -344 -134 -336
rect -119 -347 -115 -339
rect -111 -347 -107 -339
rect -103 -347 -99 -339
rect -95 -342 -91 -338
rect -87 -342 -83 -338
<< pdcontact >>
rect -176 599 -172 615
rect -168 599 -164 615
rect -160 599 -156 615
rect -146 599 -142 615
rect -138 599 -134 615
rect -130 599 -126 615
rect -121 599 -117 607
rect -113 599 -109 607
rect -103 599 -99 607
rect -95 599 -91 607
rect -87 599 -83 607
rect -79 599 -75 607
rect -176 504 -172 520
rect -168 504 -164 520
rect -160 504 -156 520
rect -146 504 -142 520
rect -138 504 -134 520
rect -130 504 -126 520
rect -121 504 -117 512
rect -113 504 -109 512
rect -103 504 -99 512
rect -95 504 -91 512
rect -87 504 -83 512
rect -79 504 -75 512
rect -175 408 -171 424
rect -167 408 -163 424
rect -159 408 -155 424
rect -145 408 -141 424
rect -137 408 -133 424
rect -129 408 -125 424
rect 32 422 36 438
rect 40 422 44 438
rect 48 422 52 438
rect 62 422 66 438
rect 70 422 74 438
rect 78 422 82 438
rect 87 422 91 430
rect 95 422 99 430
rect 105 422 109 430
rect 113 422 117 430
rect 121 422 125 430
rect 129 422 133 430
rect -120 408 -116 416
rect -112 408 -108 416
rect -102 408 -98 416
rect -94 408 -90 416
rect -86 408 -82 416
rect -78 408 -74 416
rect 155 401 159 409
rect 163 401 167 409
rect 171 401 175 409
rect 199 401 203 409
rect 207 401 211 409
rect 215 401 219 409
rect 243 401 247 409
rect 251 401 255 409
rect 259 401 263 409
rect 287 401 291 409
rect 295 401 299 409
rect 303 401 307 409
rect 331 401 335 409
rect 339 401 343 409
rect 347 401 351 409
rect -171 314 -167 330
rect -163 314 -159 330
rect -155 314 -151 330
rect -141 314 -137 330
rect -133 314 -129 330
rect -125 314 -121 330
rect 11 327 19 331
rect -116 314 -112 322
rect -108 314 -104 322
rect -98 314 -94 322
rect -90 314 -86 322
rect -82 314 -78 322
rect -74 314 -70 322
rect 11 319 19 323
rect 65 323 69 331
rect 73 323 77 331
rect 671 325 679 329
rect 11 309 19 313
rect 671 317 679 321
rect 745 312 749 328
rect 753 312 757 328
rect 761 312 765 328
rect 775 312 779 328
rect 783 312 787 328
rect 791 312 795 328
rect 800 312 804 320
rect 808 312 812 320
rect 818 312 822 320
rect 826 312 830 320
rect 834 312 838 320
rect 842 312 846 320
rect 671 307 679 311
rect 11 301 19 305
rect 671 299 679 303
rect 11 291 19 295
rect 671 289 679 293
rect 11 283 19 287
rect 671 281 679 285
rect 10 259 18 263
rect 60 259 64 267
rect 68 259 72 267
rect 10 251 18 255
rect 10 241 18 245
rect 671 250 679 254
rect 671 242 679 246
rect -170 215 -166 231
rect -162 215 -158 231
rect -154 215 -150 231
rect -140 215 -136 231
rect -132 215 -128 231
rect -124 215 -120 231
rect 10 233 18 237
rect 671 232 679 236
rect -115 215 -111 223
rect -107 215 -103 223
rect -97 215 -93 223
rect -89 215 -85 223
rect -81 215 -77 223
rect -73 215 -69 223
rect 10 223 18 227
rect 671 224 679 228
rect 10 215 18 219
rect 671 214 679 218
rect 745 217 749 233
rect 753 217 757 233
rect 761 217 765 233
rect 775 217 779 233
rect 783 217 787 233
rect 791 217 795 233
rect 800 217 804 225
rect 808 217 812 225
rect 818 217 822 225
rect 826 217 830 225
rect 834 217 838 225
rect 842 217 846 225
rect 671 206 679 210
rect 10 192 18 196
rect 60 192 64 200
rect 68 192 72 200
rect 10 184 18 188
rect 10 174 18 178
rect 207 183 211 191
rect 215 183 219 191
rect 254 183 258 191
rect 262 183 266 191
rect 288 183 292 191
rect 296 183 300 191
rect 335 183 339 191
rect 343 183 347 191
rect 369 183 373 191
rect 377 183 381 191
rect 416 183 420 191
rect 424 183 428 191
rect 450 183 454 191
rect 458 183 462 191
rect 497 183 501 191
rect 505 183 509 191
rect 531 183 535 191
rect 539 183 543 191
rect 578 183 582 191
rect 586 183 590 191
rect 10 166 18 170
rect -169 139 -165 155
rect -161 139 -157 155
rect -153 139 -149 155
rect -139 139 -135 155
rect -131 139 -127 155
rect -123 139 -119 155
rect 10 156 18 160
rect 10 148 18 152
rect 671 165 679 169
rect 671 157 679 161
rect 671 147 679 151
rect -114 139 -110 147
rect -106 139 -102 147
rect -96 139 -92 147
rect -88 139 -84 147
rect -80 139 -76 147
rect -72 139 -68 147
rect 671 139 679 143
rect 10 122 18 126
rect 60 122 64 130
rect 68 122 72 130
rect 671 129 679 133
rect 10 114 18 118
rect 10 104 18 108
rect 671 121 679 125
rect 746 121 750 137
rect 754 121 758 137
rect 762 121 766 137
rect 776 121 780 137
rect 784 121 788 137
rect 792 121 796 137
rect 801 121 805 129
rect 809 121 813 129
rect 819 121 823 129
rect 827 121 831 129
rect 835 121 839 129
rect 843 121 847 129
rect 10 96 18 100
rect 10 86 18 90
rect 10 78 18 82
rect 680 78 688 82
rect 680 70 688 74
rect 680 60 688 64
rect -174 35 -170 51
rect -166 35 -162 51
rect -158 35 -154 51
rect -144 35 -140 51
rect -136 35 -132 51
rect -128 35 -124 51
rect 10 50 18 54
rect 60 50 64 58
rect 68 50 72 58
rect 680 52 688 56
rect -119 35 -115 43
rect -111 35 -107 43
rect -101 35 -97 43
rect -93 35 -89 43
rect -85 35 -81 43
rect -77 35 -73 43
rect 10 42 18 46
rect 10 32 18 36
rect 680 42 688 46
rect 680 34 688 38
rect 10 24 18 28
rect 750 27 754 43
rect 758 27 762 43
rect 766 27 770 43
rect 780 27 784 43
rect 788 27 792 43
rect 796 27 800 43
rect 805 27 809 35
rect 813 27 817 35
rect 823 27 827 35
rect 831 27 835 35
rect 839 27 843 35
rect 847 27 851 35
rect 10 14 18 18
rect 10 6 18 10
rect 680 -58 688 -54
rect -180 -79 -176 -63
rect -172 -79 -168 -63
rect -164 -79 -160 -63
rect -150 -79 -146 -63
rect -142 -79 -138 -63
rect -134 -79 -130 -63
rect 680 -66 688 -62
rect -125 -79 -121 -71
rect -117 -79 -113 -71
rect -107 -79 -103 -71
rect -99 -79 -95 -71
rect -91 -79 -87 -71
rect -83 -79 -79 -71
rect 751 -72 755 -56
rect 759 -72 763 -56
rect 767 -72 771 -56
rect 781 -72 785 -56
rect 789 -72 793 -56
rect 797 -72 801 -56
rect 806 -72 810 -64
rect 814 -72 818 -64
rect 824 -72 828 -64
rect 832 -72 836 -64
rect 840 -72 844 -64
rect 848 -72 852 -64
rect 680 -76 688 -72
rect 680 -84 688 -80
rect 680 -94 688 -90
rect 680 -102 688 -98
rect 271 -136 275 -120
rect 279 -136 283 -120
rect 287 -136 291 -120
rect 325 -136 329 -120
rect 333 -136 337 -120
rect 341 -136 345 -120
rect 373 -136 377 -120
rect 381 -136 385 -120
rect 389 -136 393 -120
rect 421 -136 425 -120
rect 429 -136 433 -120
rect 437 -136 441 -120
rect 480 -136 484 -120
rect 488 -136 492 -120
rect 496 -136 500 -120
rect 753 -177 757 -161
rect 761 -177 765 -161
rect 769 -177 773 -161
rect 783 -177 787 -161
rect 791 -177 795 -161
rect 799 -177 803 -161
rect 808 -177 812 -169
rect 816 -177 820 -169
rect 826 -177 830 -169
rect 834 -177 838 -169
rect 842 -177 846 -169
rect 850 -177 854 -169
rect -183 -212 -179 -196
rect -175 -212 -171 -196
rect -167 -212 -163 -196
rect -153 -212 -149 -196
rect -145 -212 -141 -196
rect -137 -212 -133 -196
rect -128 -212 -124 -204
rect -120 -212 -116 -204
rect -110 -212 -106 -204
rect -102 -212 -98 -204
rect -94 -212 -90 -204
rect -86 -212 -82 -204
rect -184 -324 -180 -308
rect -176 -324 -172 -308
rect -168 -324 -164 -308
rect -154 -324 -150 -308
rect -146 -324 -142 -308
rect -138 -324 -134 -308
rect -129 -324 -125 -316
rect -121 -324 -117 -316
rect -111 -324 -107 -316
rect -103 -324 -99 -316
rect -95 -324 -91 -316
rect -87 -324 -83 -316
<< polysilicon >>
rect -171 615 -169 618
rect -163 615 -161 624
rect -141 615 -139 618
rect -133 615 -131 627
rect -116 607 -114 620
rect -98 607 -96 613
rect -82 607 -80 613
rect -171 585 -169 599
rect -163 591 -161 599
rect -141 587 -139 599
rect -133 587 -131 599
rect -116 593 -114 599
rect -98 592 -96 599
rect -106 590 -96 592
rect -171 578 -169 581
rect -106 584 -104 590
rect -98 584 -96 587
rect -82 585 -80 599
rect -141 568 -139 579
rect -133 576 -131 579
rect -82 577 -80 581
rect -106 573 -104 576
rect -98 573 -96 576
rect -171 520 -169 523
rect -163 520 -161 529
rect -141 520 -139 523
rect -133 520 -131 532
rect -116 512 -114 525
rect -98 512 -96 518
rect -82 512 -80 518
rect -171 490 -169 504
rect -163 496 -161 504
rect -141 492 -139 504
rect -133 492 -131 504
rect -116 498 -114 504
rect -98 497 -96 504
rect -106 495 -96 497
rect -171 483 -169 486
rect -106 489 -104 495
rect -98 489 -96 492
rect -82 490 -80 504
rect -141 473 -139 484
rect -133 481 -131 484
rect -82 482 -80 486
rect -106 478 -104 481
rect -98 478 -96 481
rect 37 438 39 441
rect 45 438 47 447
rect 67 438 69 441
rect 75 438 77 450
rect -170 424 -168 427
rect -162 424 -160 433
rect -140 424 -138 427
rect -132 424 -130 436
rect -115 416 -113 429
rect 92 430 94 443
rect 110 430 112 436
rect 126 430 128 436
rect -97 416 -95 422
rect -81 416 -79 422
rect 37 408 39 422
rect 45 414 47 422
rect 67 410 69 422
rect 75 410 77 422
rect 92 416 94 422
rect 110 415 112 422
rect 102 413 112 415
rect -170 394 -168 408
rect -162 400 -160 408
rect -140 396 -138 408
rect -132 396 -130 408
rect -115 402 -113 408
rect -97 401 -95 408
rect -105 399 -95 401
rect -170 387 -168 390
rect -105 393 -103 399
rect -97 393 -95 396
rect -81 394 -79 408
rect 37 401 39 404
rect 102 407 104 413
rect 110 407 112 410
rect 126 408 128 422
rect 160 409 162 423
rect 168 409 170 423
rect 204 409 206 423
rect 212 409 214 423
rect 248 409 250 423
rect 256 409 258 423
rect 292 409 294 423
rect 300 409 302 423
rect 336 409 338 423
rect 344 409 346 423
rect -140 377 -138 388
rect -132 385 -130 388
rect 67 391 69 402
rect 75 399 77 402
rect 126 400 128 404
rect 102 396 104 399
rect 110 396 112 399
rect -81 386 -79 390
rect -105 382 -103 385
rect -97 382 -95 385
rect 160 383 162 401
rect 168 383 170 401
rect 204 383 206 401
rect 212 383 214 401
rect 248 383 250 401
rect 256 383 258 401
rect 292 383 294 401
rect 300 383 302 401
rect 336 383 338 401
rect 344 383 346 401
rect 160 371 162 375
rect 168 371 170 375
rect 204 371 206 375
rect 212 371 214 375
rect 248 371 250 375
rect 256 371 258 375
rect 292 371 294 375
rect 300 371 302 375
rect 336 371 338 375
rect 344 371 346 375
rect -166 330 -164 333
rect -158 330 -156 339
rect -136 330 -134 333
rect -128 330 -126 342
rect -111 322 -109 335
rect 70 331 72 335
rect -93 322 -91 328
rect -77 322 -75 328
rect 1 324 11 326
rect 19 324 25 326
rect 28 324 31 326
rect 35 324 44 326
rect 750 328 752 331
rect 758 328 760 337
rect 780 328 782 331
rect 788 328 790 340
rect -166 300 -164 314
rect -158 306 -156 314
rect -136 302 -134 314
rect -128 302 -126 314
rect -111 308 -109 314
rect -93 307 -91 314
rect -101 305 -91 307
rect -166 293 -164 296
rect -101 299 -99 305
rect -93 299 -91 302
rect -77 300 -75 314
rect 7 306 11 308
rect 19 306 31 308
rect 35 306 38 308
rect 70 306 72 323
rect 661 322 671 324
rect 679 322 685 324
rect 688 322 691 324
rect 695 322 704 324
rect 805 320 807 333
rect 823 320 825 326
rect 839 320 841 326
rect 667 304 671 306
rect 679 304 691 306
rect 695 304 698 306
rect -136 283 -134 294
rect -128 291 -126 294
rect 70 299 72 302
rect 750 298 752 312
rect 758 304 760 312
rect 780 300 782 312
rect 788 300 790 312
rect 805 306 807 312
rect 823 305 825 312
rect 815 303 825 305
rect -77 292 -75 296
rect -101 288 -99 291
rect -93 288 -91 291
rect 3 288 11 290
rect 19 288 35 290
rect 39 288 42 290
rect 750 291 752 294
rect 815 297 817 303
rect 823 297 825 300
rect 839 298 841 312
rect 663 286 671 288
rect 679 286 695 288
rect 699 286 702 288
rect 780 281 782 292
rect 788 289 790 292
rect 839 290 841 294
rect 815 286 817 289
rect 823 286 825 289
rect 65 267 67 271
rect 0 256 10 258
rect 18 256 24 258
rect 27 256 30 258
rect 34 256 43 258
rect -165 231 -163 234
rect -157 231 -155 240
rect -135 231 -133 234
rect -127 231 -125 243
rect 65 242 67 259
rect 661 247 671 249
rect 679 247 685 249
rect 688 247 691 249
rect 695 247 704 249
rect 6 238 10 240
rect 18 238 30 240
rect 34 238 37 240
rect -110 223 -108 236
rect 65 235 67 238
rect 750 233 752 236
rect 758 233 760 242
rect 780 233 782 236
rect 788 233 790 245
rect 667 229 671 231
rect 679 229 691 231
rect 695 229 698 231
rect -92 223 -90 229
rect -76 223 -74 229
rect 2 220 10 222
rect 18 220 34 222
rect 38 220 41 222
rect -165 201 -163 215
rect -157 207 -155 215
rect -135 203 -133 215
rect -127 203 -125 215
rect -110 209 -108 215
rect -92 208 -90 215
rect -100 206 -90 208
rect -165 194 -163 197
rect -100 200 -98 206
rect -92 200 -90 203
rect -76 201 -74 215
rect 805 225 807 238
rect 823 225 825 231
rect 839 225 841 231
rect 663 211 671 213
rect 679 211 695 213
rect 699 211 702 213
rect -135 184 -133 195
rect -127 192 -125 195
rect 65 200 67 204
rect 750 203 752 217
rect 758 209 760 217
rect 780 205 782 217
rect 788 205 790 217
rect 805 211 807 217
rect 823 210 825 217
rect 815 208 825 210
rect -76 193 -74 197
rect -100 189 -98 192
rect -92 189 -90 192
rect 0 189 10 191
rect 18 189 24 191
rect 27 189 30 191
rect 34 189 43 191
rect 65 175 67 192
rect 212 191 214 199
rect 259 191 261 199
rect 293 191 295 199
rect 340 191 342 199
rect 374 191 376 199
rect 421 191 423 199
rect 455 191 457 199
rect 502 191 504 199
rect 536 191 538 199
rect 583 191 585 199
rect 750 196 752 199
rect 815 202 817 208
rect 823 202 825 205
rect 839 203 841 217
rect 780 186 782 197
rect 788 194 790 197
rect 839 195 841 199
rect 815 191 817 194
rect 823 191 825 194
rect 6 171 10 173
rect 18 171 30 173
rect 34 171 37 173
rect 212 174 214 183
rect 259 174 261 183
rect 293 174 295 183
rect 340 174 342 183
rect 374 174 376 183
rect 421 174 423 183
rect 455 174 457 183
rect 502 174 504 183
rect 536 174 538 183
rect 583 174 585 183
rect -164 155 -162 158
rect -156 155 -154 164
rect -134 155 -132 158
rect -126 155 -124 167
rect 65 168 67 171
rect 212 166 214 169
rect 259 165 261 168
rect 293 166 295 169
rect -109 147 -107 160
rect 2 153 10 155
rect 18 153 34 155
rect 38 153 41 155
rect -91 147 -89 153
rect -75 147 -73 153
rect 212 152 214 162
rect 340 165 342 168
rect 374 166 376 169
rect 259 152 261 161
rect 293 152 295 162
rect 421 165 423 168
rect 455 166 457 169
rect 340 152 342 161
rect 374 152 376 162
rect 502 165 504 168
rect 536 166 538 169
rect 421 152 423 161
rect 455 152 457 162
rect 583 165 585 168
rect 502 152 504 161
rect 536 152 538 162
rect 661 162 671 164
rect 679 162 685 164
rect 688 162 691 164
rect 695 162 704 164
rect 583 152 585 161
rect 667 144 671 146
rect 679 144 691 146
rect 695 144 698 146
rect -164 125 -162 139
rect -156 131 -154 139
rect -134 127 -132 139
rect -126 127 -124 139
rect -109 133 -107 139
rect -91 132 -89 139
rect -99 130 -89 132
rect -164 118 -162 121
rect -99 124 -97 130
rect -91 124 -89 127
rect -75 125 -73 139
rect 751 137 753 140
rect 759 137 761 146
rect 781 137 783 140
rect 789 137 791 149
rect 65 130 67 134
rect -134 108 -132 119
rect -126 116 -124 119
rect 663 126 671 128
rect 679 126 695 128
rect 699 126 702 128
rect -75 117 -73 121
rect 0 119 10 121
rect 18 119 24 121
rect 27 119 30 121
rect 34 119 43 121
rect -99 113 -97 116
rect -91 113 -89 116
rect 65 105 67 122
rect 806 129 808 142
rect 824 129 826 135
rect 840 129 842 135
rect 751 107 753 121
rect 759 113 761 121
rect 781 109 783 121
rect 789 109 791 121
rect 806 115 808 121
rect 824 114 826 121
rect 816 112 826 114
rect 6 101 10 103
rect 18 101 30 103
rect 34 101 37 103
rect 65 98 67 101
rect 751 100 753 103
rect 816 106 818 112
rect 824 106 826 109
rect 840 107 842 121
rect 781 90 783 101
rect 789 98 791 101
rect 840 99 842 103
rect 816 95 818 98
rect 824 95 826 98
rect 2 83 10 85
rect 18 83 34 85
rect 38 83 41 85
rect 670 75 680 77
rect 688 75 694 77
rect 697 75 700 77
rect 704 75 713 77
rect -169 51 -167 54
rect -161 51 -159 60
rect -139 51 -137 54
rect -131 51 -129 63
rect 65 58 67 62
rect -114 43 -112 56
rect 676 57 680 59
rect 688 57 700 59
rect 704 57 707 59
rect -96 43 -94 49
rect -80 43 -78 49
rect 0 47 10 49
rect 18 47 24 49
rect 27 47 30 49
rect 34 47 43 49
rect -169 21 -167 35
rect -161 27 -159 35
rect -139 23 -137 35
rect -131 23 -129 35
rect -114 29 -112 35
rect -96 28 -94 35
rect -104 26 -94 28
rect -169 14 -167 17
rect -104 20 -102 26
rect -96 20 -94 23
rect -80 21 -78 35
rect 65 33 67 50
rect 755 43 757 46
rect 763 43 765 52
rect 785 43 787 46
rect 793 43 795 55
rect 672 39 680 41
rect 688 39 704 41
rect 708 39 711 41
rect 6 29 10 31
rect 18 29 30 31
rect 34 29 37 31
rect 65 26 67 29
rect 810 35 812 48
rect 828 35 830 41
rect 844 35 846 41
rect -139 4 -137 15
rect -131 12 -129 15
rect -80 13 -78 17
rect 755 13 757 27
rect 763 19 765 27
rect 785 15 787 27
rect 793 15 795 27
rect 810 21 812 27
rect 828 20 830 27
rect 820 18 830 20
rect -104 9 -102 12
rect -96 9 -94 12
rect 2 11 10 13
rect 18 11 34 13
rect 38 11 41 13
rect 755 6 757 9
rect 820 12 822 18
rect 828 12 830 15
rect 844 13 846 27
rect 785 -4 787 7
rect 793 4 795 7
rect 844 5 846 9
rect 820 1 822 4
rect 828 1 830 4
rect -175 -63 -173 -60
rect -167 -63 -165 -54
rect -145 -63 -143 -60
rect -137 -63 -135 -51
rect -120 -71 -118 -58
rect 756 -56 758 -53
rect 764 -56 766 -47
rect 786 -56 788 -53
rect 794 -56 796 -44
rect 670 -61 680 -59
rect 688 -61 694 -59
rect 697 -61 700 -59
rect 704 -61 713 -59
rect -102 -71 -100 -65
rect -86 -71 -84 -65
rect 811 -64 813 -51
rect 829 -64 831 -58
rect 845 -64 847 -58
rect 676 -79 680 -77
rect 688 -79 700 -77
rect 704 -79 707 -77
rect -175 -93 -173 -79
rect -167 -87 -165 -79
rect -145 -91 -143 -79
rect -137 -91 -135 -79
rect -120 -85 -118 -79
rect -102 -86 -100 -79
rect -110 -88 -100 -86
rect -175 -100 -173 -97
rect -110 -94 -108 -88
rect -102 -94 -100 -91
rect -86 -93 -84 -79
rect 756 -86 758 -72
rect 764 -80 766 -72
rect 786 -84 788 -72
rect 794 -84 796 -72
rect 811 -78 813 -72
rect 829 -79 831 -72
rect 821 -81 831 -79
rect -145 -110 -143 -99
rect -137 -102 -135 -99
rect 756 -93 758 -90
rect 821 -87 823 -81
rect 829 -87 831 -84
rect 845 -86 847 -72
rect 672 -97 680 -95
rect 688 -97 704 -95
rect 708 -97 711 -95
rect -86 -101 -84 -97
rect 276 -100 278 -97
rect 284 -100 286 -97
rect 330 -100 332 -97
rect 338 -100 340 -97
rect 378 -100 380 -97
rect 386 -100 388 -97
rect 426 -100 428 -97
rect 434 -100 436 -97
rect 485 -100 487 -97
rect 493 -100 495 -97
rect -110 -105 -108 -102
rect -102 -105 -100 -102
rect 786 -103 788 -92
rect 794 -95 796 -92
rect 845 -94 847 -90
rect 821 -98 823 -95
rect 829 -98 831 -95
rect 276 -120 278 -104
rect 284 -120 286 -104
rect 330 -120 332 -104
rect 338 -120 340 -104
rect 378 -120 380 -104
rect 386 -120 388 -104
rect 426 -120 428 -104
rect 434 -120 436 -104
rect 485 -120 487 -104
rect 493 -120 495 -104
rect 276 -147 278 -136
rect 284 -147 286 -136
rect 330 -147 332 -136
rect 338 -147 340 -136
rect 378 -147 380 -136
rect 386 -147 388 -136
rect 426 -147 428 -136
rect 434 -147 436 -136
rect 485 -147 487 -136
rect 493 -147 495 -136
rect 758 -161 760 -158
rect 766 -161 768 -152
rect 788 -161 790 -158
rect 796 -161 798 -149
rect 813 -169 815 -156
rect 831 -169 833 -163
rect 847 -169 849 -163
rect -178 -196 -176 -193
rect -170 -196 -168 -187
rect -148 -196 -146 -193
rect -140 -196 -138 -184
rect 758 -191 760 -177
rect 766 -185 768 -177
rect 788 -189 790 -177
rect 796 -189 798 -177
rect 813 -183 815 -177
rect 831 -184 833 -177
rect 823 -186 833 -184
rect -123 -204 -121 -191
rect 758 -198 760 -195
rect 823 -192 825 -186
rect 831 -192 833 -189
rect 847 -191 849 -177
rect -105 -204 -103 -198
rect -89 -204 -87 -198
rect 788 -208 790 -197
rect 796 -200 798 -197
rect 847 -199 849 -195
rect 823 -203 825 -200
rect 831 -203 833 -200
rect -178 -226 -176 -212
rect -170 -220 -168 -212
rect -148 -224 -146 -212
rect -140 -224 -138 -212
rect -123 -218 -121 -212
rect -105 -219 -103 -212
rect -113 -221 -103 -219
rect -178 -233 -176 -230
rect -113 -227 -111 -221
rect -105 -227 -103 -224
rect -89 -226 -87 -212
rect -148 -243 -146 -232
rect -140 -235 -138 -232
rect -89 -234 -87 -230
rect -113 -238 -111 -235
rect -105 -238 -103 -235
rect -179 -308 -177 -305
rect -171 -308 -169 -299
rect -149 -308 -147 -305
rect -141 -308 -139 -296
rect -124 -316 -122 -303
rect -106 -316 -104 -310
rect -90 -316 -88 -310
rect -179 -338 -177 -324
rect -171 -332 -169 -324
rect -149 -336 -147 -324
rect -141 -336 -139 -324
rect -124 -330 -122 -324
rect -106 -331 -104 -324
rect -114 -333 -104 -331
rect -179 -345 -177 -342
rect -114 -339 -112 -333
rect -106 -339 -104 -336
rect -90 -338 -88 -324
rect -149 -355 -147 -344
rect -141 -347 -139 -344
rect -90 -346 -88 -342
rect -114 -350 -112 -347
rect -106 -350 -104 -347
<< polycontact >>
rect -164 624 -160 628
rect -137 623 -133 627
rect -114 616 -110 620
rect -175 588 -171 592
rect -110 588 -106 592
rect -86 588 -82 592
rect -99 569 -95 573
rect -142 564 -138 568
rect -164 529 -160 533
rect -137 528 -133 532
rect -114 521 -110 525
rect -175 493 -171 497
rect -110 493 -106 497
rect -86 493 -82 497
rect -99 474 -95 478
rect -142 469 -138 473
rect 44 447 48 451
rect 71 446 75 450
rect -163 433 -159 437
rect -136 432 -132 436
rect -113 425 -109 429
rect 94 439 98 443
rect 159 423 163 427
rect 167 423 171 427
rect 203 423 207 427
rect 211 423 215 427
rect 247 423 251 427
rect 255 423 259 427
rect 291 423 295 427
rect 299 423 303 427
rect 335 423 339 427
rect 343 423 347 427
rect 33 411 37 415
rect 98 411 102 415
rect -174 397 -170 401
rect -109 397 -105 401
rect -85 397 -81 401
rect 122 411 126 415
rect 109 392 113 396
rect 66 387 70 391
rect -98 378 -94 382
rect -141 373 -137 377
rect -159 339 -155 343
rect -132 338 -128 342
rect 757 337 761 341
rect -109 331 -105 335
rect 1 320 5 324
rect 40 320 44 324
rect 784 336 788 340
rect -170 303 -166 307
rect -105 303 -101 307
rect -81 303 -77 307
rect 65 313 70 319
rect 661 318 665 322
rect 700 318 704 322
rect 807 329 811 333
rect 22 302 26 306
rect 682 300 686 304
rect 746 301 750 305
rect 811 301 815 305
rect 3 290 7 294
rect 663 288 667 292
rect 835 301 839 305
rect -94 284 -90 288
rect -137 279 -133 283
rect 822 282 826 286
rect 779 277 783 281
rect 0 252 4 256
rect 39 252 43 256
rect 60 245 65 251
rect -158 240 -154 244
rect -131 239 -127 243
rect 661 243 665 247
rect 700 243 704 247
rect 757 242 761 246
rect -108 232 -104 236
rect 21 234 25 238
rect 784 241 788 245
rect 2 222 6 226
rect 682 225 686 229
rect -169 204 -165 208
rect -104 204 -100 208
rect -80 204 -76 208
rect 663 213 667 217
rect 807 234 811 238
rect 746 206 750 210
rect 811 206 815 210
rect -93 185 -89 189
rect 0 185 4 189
rect 39 185 43 189
rect -136 180 -132 184
rect 60 178 65 184
rect 214 194 218 198
rect 261 194 265 198
rect 295 194 299 198
rect 342 194 346 198
rect 376 194 380 198
rect 423 194 427 198
rect 457 194 461 198
rect 504 194 508 198
rect 538 194 542 198
rect 585 194 589 198
rect 835 206 839 210
rect 822 187 826 191
rect 779 182 783 186
rect -157 164 -153 168
rect -130 163 -126 167
rect 21 167 25 171
rect -107 156 -103 160
rect 2 155 6 159
rect 214 154 218 158
rect 261 154 265 158
rect 295 154 299 158
rect 342 154 346 158
rect 376 154 380 158
rect 423 154 427 158
rect 457 154 461 158
rect 504 154 508 158
rect 538 154 542 158
rect 661 158 665 162
rect 585 154 589 158
rect 700 158 704 162
rect 758 146 762 150
rect 682 140 686 144
rect -168 128 -164 132
rect -103 128 -99 132
rect -79 128 -75 132
rect 785 145 789 149
rect 663 128 667 132
rect 0 115 4 119
rect 39 115 43 119
rect -92 109 -88 113
rect 60 108 65 114
rect -135 104 -131 108
rect 808 138 812 142
rect 747 110 751 114
rect 812 110 816 114
rect 21 97 25 101
rect 836 110 840 114
rect 823 91 827 95
rect 2 85 6 89
rect 780 86 784 90
rect 670 71 674 75
rect 709 71 713 75
rect -162 60 -158 64
rect -135 59 -131 63
rect -112 52 -108 56
rect 691 53 695 57
rect 762 52 766 56
rect 0 43 4 47
rect 39 43 43 47
rect 60 36 65 42
rect -173 24 -169 28
rect -108 24 -104 28
rect -84 24 -80 28
rect 672 41 676 45
rect 789 51 793 55
rect 21 25 25 29
rect 812 44 816 48
rect 2 13 6 17
rect 751 16 755 20
rect 816 16 820 20
rect -97 5 -93 9
rect 840 16 844 20
rect -140 0 -136 4
rect 827 -3 831 1
rect 784 -8 788 -4
rect 763 -47 767 -43
rect -168 -54 -164 -50
rect -141 -55 -137 -51
rect -118 -62 -114 -58
rect 790 -48 794 -44
rect 670 -65 674 -61
rect 709 -65 713 -61
rect 813 -55 817 -51
rect -179 -90 -175 -86
rect -114 -90 -110 -86
rect -90 -90 -86 -86
rect 691 -83 695 -79
rect 752 -83 756 -79
rect 817 -83 821 -79
rect 672 -95 676 -91
rect 841 -83 845 -79
rect 828 -102 832 -98
rect -103 -109 -99 -105
rect -146 -114 -142 -110
rect 785 -107 789 -103
rect 275 -151 279 -147
rect 283 -151 287 -147
rect 329 -151 333 -147
rect 337 -151 341 -147
rect 377 -151 381 -147
rect 385 -151 389 -147
rect 425 -151 429 -147
rect 433 -151 437 -147
rect 484 -151 488 -147
rect 492 -151 496 -147
rect 765 -152 769 -148
rect 792 -153 796 -149
rect 815 -160 819 -156
rect -171 -187 -167 -183
rect -144 -188 -140 -184
rect 754 -188 758 -184
rect 819 -188 823 -184
rect -121 -195 -117 -191
rect 843 -188 847 -184
rect 830 -207 834 -203
rect 787 -212 791 -208
rect -182 -223 -178 -219
rect -117 -223 -113 -219
rect -93 -223 -89 -219
rect -106 -242 -102 -238
rect -149 -247 -145 -243
rect -172 -299 -168 -295
rect -145 -300 -141 -296
rect -122 -307 -118 -303
rect -183 -335 -179 -331
rect -118 -335 -114 -331
rect -94 -335 -90 -331
rect -107 -354 -103 -350
rect -150 -359 -146 -355
<< metal1 >>
rect -164 628 -160 631
rect -176 615 -172 624
rect -153 623 -137 627
rect -182 588 -175 592
rect -160 589 -156 599
rect -153 589 -149 623
rect -146 615 -142 620
rect -110 616 -107 620
rect -121 607 -117 616
rect -103 607 -99 613
rect -87 607 -83 613
rect -168 586 -149 589
rect -130 592 -126 599
rect -113 592 -109 599
rect -95 592 -91 599
rect -79 592 -75 599
rect -72 592 -58 593
rect -130 588 -110 592
rect -95 588 -86 592
rect -79 588 -58 592
rect -130 587 -126 588
rect -168 585 -164 586
rect -176 578 -172 581
rect -95 584 -91 588
rect -79 585 -75 588
rect -146 577 -142 579
rect -150 573 -142 577
rect -87 576 -83 581
rect -111 572 -107 576
rect -99 566 -95 569
rect -142 561 -138 564
rect -63 561 -58 588
rect -63 556 -8 561
rect -164 533 -160 536
rect -176 520 -172 529
rect -153 528 -137 532
rect -182 493 -175 497
rect -160 494 -156 504
rect -153 494 -149 528
rect -146 520 -142 525
rect -110 521 -107 525
rect -121 512 -117 521
rect -103 512 -99 518
rect -87 512 -83 518
rect -168 491 -149 494
rect -130 497 -126 504
rect -113 497 -109 504
rect -95 497 -91 504
rect -79 497 -75 504
rect -72 497 -19 498
rect -130 493 -110 497
rect -95 493 -86 497
rect -79 493 -19 497
rect -130 492 -126 493
rect -168 490 -164 491
rect -176 483 -172 486
rect -95 489 -91 493
rect -79 490 -75 493
rect -146 482 -142 484
rect -150 478 -142 482
rect -87 481 -83 486
rect -111 477 -107 481
rect -99 471 -95 474
rect -142 466 -138 469
rect -163 437 -159 440
rect -175 424 -171 433
rect -152 432 -136 436
rect -181 397 -174 401
rect -159 398 -155 408
rect -152 398 -148 432
rect -145 424 -141 429
rect -109 425 -106 429
rect -120 416 -116 425
rect -102 416 -98 422
rect -86 416 -82 422
rect -167 395 -148 398
rect -129 401 -125 408
rect -112 401 -108 408
rect -94 401 -90 408
rect -78 401 -74 408
rect -69 401 -30 402
rect -129 397 -109 401
rect -94 397 -85 401
rect -78 397 -30 401
rect -129 396 -125 397
rect -167 394 -163 395
rect -175 387 -171 390
rect -94 393 -90 397
rect -78 394 -74 397
rect -145 386 -141 388
rect -149 382 -141 386
rect -86 385 -82 390
rect -110 381 -106 385
rect -98 375 -94 378
rect -141 370 -137 373
rect -159 343 -155 346
rect -171 330 -167 339
rect -148 338 -132 342
rect -177 303 -170 307
rect -155 304 -151 314
rect -148 304 -144 338
rect -141 330 -137 335
rect -105 331 -102 335
rect -116 322 -112 331
rect -98 322 -94 328
rect -82 322 -78 328
rect -163 301 -144 304
rect -125 307 -121 314
rect -108 307 -104 314
rect -90 307 -86 314
rect -74 307 -70 314
rect -64 307 -40 308
rect -125 303 -105 307
rect -90 303 -81 307
rect -74 303 -40 307
rect -125 302 -121 303
rect -163 300 -159 301
rect -171 293 -167 296
rect -90 299 -86 303
rect -74 300 -70 303
rect -141 292 -137 294
rect -145 288 -137 292
rect -82 291 -78 296
rect -106 287 -102 291
rect -94 281 -90 284
rect -137 276 -133 279
rect -158 244 -154 247
rect -170 231 -166 240
rect -147 239 -131 243
rect -176 204 -169 208
rect -154 205 -150 215
rect -147 205 -143 239
rect -140 231 -136 236
rect -104 232 -101 236
rect -115 223 -111 232
rect -97 223 -93 229
rect -81 223 -77 229
rect -162 202 -143 205
rect -124 208 -120 215
rect -107 208 -103 215
rect -89 208 -85 215
rect -73 208 -69 215
rect -64 208 -49 209
rect -124 204 -104 208
rect -89 204 -80 208
rect -73 204 -49 208
rect -124 203 -120 204
rect -162 201 -158 202
rect -170 194 -166 197
rect -89 200 -85 204
rect -73 201 -69 204
rect -140 193 -136 195
rect -144 189 -136 193
rect -81 192 -77 197
rect -105 188 -101 192
rect -93 182 -89 185
rect -136 177 -132 180
rect -157 168 -153 171
rect -169 155 -165 164
rect -146 163 -130 167
rect -175 128 -168 132
rect -153 129 -149 139
rect -146 129 -142 163
rect -139 155 -135 160
rect -103 156 -100 160
rect -114 147 -110 156
rect -96 147 -92 153
rect -80 147 -76 153
rect -161 126 -142 129
rect -123 132 -119 139
rect -106 132 -102 139
rect -88 132 -84 139
rect -72 132 -68 139
rect -54 141 -49 204
rect -45 153 -40 303
rect -35 178 -30 397
rect -24 240 -19 493
rect -13 311 -8 556
rect 44 451 48 454
rect 32 438 36 447
rect 55 446 71 450
rect 26 411 33 415
rect 48 412 52 422
rect 55 412 59 446
rect 62 438 66 443
rect 98 439 101 443
rect 87 430 91 439
rect 105 430 109 436
rect 121 430 125 436
rect 159 427 163 430
rect 167 427 171 430
rect 203 427 207 430
rect 211 427 215 430
rect 247 427 251 430
rect 255 427 259 430
rect 291 427 295 430
rect 299 427 303 430
rect 335 427 339 430
rect 343 427 347 430
rect 40 409 59 412
rect 78 415 82 422
rect 95 415 99 422
rect 113 415 117 422
rect 129 415 133 422
rect 155 415 175 419
rect 78 411 98 415
rect 113 411 122 415
rect 129 411 142 415
rect 78 410 82 411
rect 40 408 44 409
rect 32 401 36 404
rect 113 407 117 411
rect 129 408 133 411
rect 62 400 66 402
rect 58 396 66 400
rect 121 399 125 404
rect 97 395 101 399
rect 109 389 113 392
rect 136 393 142 411
rect 155 409 159 415
rect 171 409 175 415
rect 199 415 219 419
rect 199 409 203 415
rect 215 409 219 415
rect 243 415 263 419
rect 243 409 247 415
rect 259 409 263 415
rect 287 415 307 419
rect 287 409 291 415
rect 303 409 307 415
rect 331 415 351 419
rect 331 409 335 415
rect 347 409 351 415
rect 136 387 144 393
rect 163 392 167 401
rect 207 392 211 401
rect 163 387 189 392
rect 207 387 224 392
rect 66 384 70 387
rect 171 383 175 387
rect 155 371 159 375
rect 184 353 189 387
rect 215 383 219 387
rect 251 392 255 401
rect 295 392 299 401
rect 307 392 313 397
rect 339 392 343 401
rect 251 387 272 392
rect 295 387 319 392
rect 339 387 606 392
rect 259 383 263 387
rect 199 371 203 375
rect 243 371 247 375
rect 184 348 246 353
rect 65 331 69 337
rect 19 327 31 331
rect 1 311 5 320
rect 19 319 31 323
rect -13 306 5 311
rect 19 309 31 313
rect 1 305 5 306
rect 1 301 11 305
rect 40 305 44 320
rect 57 313 65 319
rect 73 315 77 323
rect 96 315 102 326
rect 73 309 102 315
rect 73 306 77 309
rect 3 294 7 301
rect 22 300 26 302
rect 35 301 44 305
rect 40 295 44 301
rect 65 297 69 302
rect 19 291 35 295
rect 39 291 44 295
rect 3 283 11 287
rect 39 283 44 287
rect 267 284 272 387
rect 303 383 318 387
rect 347 383 351 387
rect 287 371 291 375
rect 307 308 318 383
rect 331 371 335 375
rect 307 303 523 308
rect 307 284 313 303
rect 267 279 436 284
rect 26 272 30 279
rect 23 266 30 272
rect 60 267 64 273
rect 26 263 29 266
rect 18 259 30 263
rect 0 240 4 252
rect 18 251 30 255
rect 18 241 30 245
rect -24 237 4 240
rect -24 235 10 237
rect 0 233 10 235
rect 39 237 43 252
rect 53 245 60 251
rect 68 250 72 259
rect 307 250 313 279
rect 68 246 313 250
rect 68 242 72 246
rect 2 226 6 233
rect 21 232 25 234
rect 34 233 43 237
rect 60 233 64 238
rect 68 237 72 238
rect 68 233 77 237
rect 39 227 43 233
rect 18 223 34 227
rect 38 223 43 227
rect 307 226 313 246
rect 518 244 523 303
rect 185 222 396 226
rect 2 215 10 219
rect 38 215 43 219
rect 8 200 29 207
rect 26 196 29 200
rect 60 200 64 206
rect 18 192 30 196
rect 185 195 189 222
rect 307 206 313 222
rect 200 202 226 206
rect 247 202 273 206
rect 281 202 313 206
rect 328 202 354 206
rect 362 202 388 206
rect 0 178 4 185
rect 18 184 30 188
rect -35 173 4 178
rect 18 174 30 178
rect 0 170 4 173
rect 0 166 10 170
rect 39 170 43 185
rect 54 178 60 184
rect 68 182 72 192
rect 167 191 189 195
rect 207 191 211 202
rect 218 194 231 198
rect 254 191 258 202
rect 265 194 275 198
rect 288 191 292 202
rect 307 198 313 202
rect 299 194 313 198
rect 167 182 171 191
rect 68 178 171 182
rect 68 175 72 178
rect 2 159 6 166
rect 21 165 25 167
rect 34 166 43 170
rect 60 166 64 171
rect 68 170 72 171
rect 68 166 77 170
rect 207 173 211 183
rect 202 169 211 173
rect 207 166 211 169
rect 39 160 43 166
rect 18 156 34 160
rect 38 156 43 160
rect 215 173 219 183
rect 262 173 266 183
rect 288 173 292 183
rect 215 169 292 173
rect 215 166 219 169
rect 262 165 266 169
rect -45 148 -23 153
rect 2 148 10 152
rect 38 148 43 152
rect 207 150 211 162
rect 288 166 292 169
rect 296 173 300 183
rect 307 173 313 194
rect 335 191 339 202
rect 346 194 355 198
rect 369 191 373 202
rect 392 198 396 222
rect 409 202 435 206
rect 443 202 469 206
rect 490 202 516 206
rect 524 202 550 206
rect 571 202 597 206
rect 380 194 396 198
rect 416 191 420 202
rect 427 194 437 198
rect 450 191 454 202
rect 461 194 483 198
rect 497 191 501 202
rect 508 194 518 198
rect 531 191 535 202
rect 542 194 560 198
rect 578 191 582 202
rect 601 198 606 387
rect 757 341 761 344
rect 687 329 690 333
rect 679 325 691 329
rect 745 328 749 337
rect 768 336 784 340
rect 661 303 665 318
rect 679 317 691 321
rect 679 307 691 311
rect 661 300 671 303
rect 650 299 671 300
rect 700 303 704 318
rect 650 294 667 299
rect 682 298 686 300
rect 695 299 704 303
rect 744 301 746 305
rect 761 302 765 312
rect 768 302 772 336
rect 775 328 779 333
rect 811 329 814 333
rect 800 320 804 329
rect 818 320 822 326
rect 834 320 838 326
rect 663 292 667 294
rect 700 293 704 299
rect 753 299 772 302
rect 791 305 795 312
rect 808 305 812 312
rect 826 305 830 312
rect 842 305 846 312
rect 791 301 811 305
rect 826 301 835 305
rect 842 301 853 305
rect 791 300 795 301
rect 753 298 757 299
rect 679 289 695 293
rect 699 289 704 293
rect 745 291 749 294
rect 826 297 830 301
rect 842 298 846 301
rect 775 290 779 292
rect 771 286 779 290
rect 834 289 838 294
rect 810 285 814 289
rect 663 281 671 285
rect 699 281 704 285
rect 822 279 826 282
rect 779 274 783 277
rect 687 254 690 258
rect 679 250 691 254
rect 661 228 665 243
rect 679 242 691 246
rect 679 232 691 236
rect 661 224 671 228
rect 700 228 704 243
rect 757 246 761 249
rect 635 218 667 224
rect 682 223 686 225
rect 695 224 704 228
rect 700 218 704 224
rect 663 217 667 218
rect 679 214 695 218
rect 699 214 704 218
rect 745 233 749 242
rect 768 241 784 245
rect 663 206 671 210
rect 699 206 704 210
rect 743 206 746 210
rect 761 207 765 217
rect 768 207 772 241
rect 775 233 779 238
rect 811 234 814 238
rect 800 225 804 234
rect 818 225 822 231
rect 834 225 838 231
rect 753 204 772 207
rect 791 210 795 217
rect 808 210 812 217
rect 826 210 830 217
rect 842 210 846 217
rect 791 206 811 210
rect 826 206 835 210
rect 842 206 853 210
rect 791 205 795 206
rect 753 203 757 204
rect 589 194 606 198
rect 745 196 749 199
rect 826 202 830 206
rect 842 203 846 206
rect 775 195 779 197
rect 771 191 779 195
rect 834 194 838 199
rect 343 173 347 183
rect 369 173 373 183
rect 296 169 373 173
rect 296 166 300 169
rect 218 154 231 158
rect 254 150 258 161
rect 265 154 276 158
rect 288 150 292 162
rect 307 159 313 169
rect 343 165 347 169
rect 369 166 373 169
rect 377 173 381 183
rect 424 173 428 183
rect 450 173 454 183
rect 377 169 454 173
rect 377 166 381 169
rect 424 165 428 169
rect 307 158 311 159
rect 299 154 311 158
rect 307 153 311 154
rect 307 150 313 153
rect 335 150 339 161
rect 346 154 358 158
rect 369 150 373 162
rect 450 166 454 169
rect 458 173 462 183
rect 505 173 509 183
rect 531 173 535 183
rect 458 169 535 173
rect 458 166 462 169
rect 505 165 509 169
rect 380 154 389 158
rect 416 150 420 161
rect 427 154 438 158
rect 450 150 454 162
rect 531 166 535 169
rect 810 190 814 194
rect 539 173 543 183
rect 586 173 590 183
rect 822 184 826 187
rect 779 179 783 182
rect 539 169 597 173
rect 539 166 543 169
rect 586 165 590 169
rect 687 169 690 173
rect 679 165 691 169
rect 461 154 470 158
rect 497 150 501 161
rect 508 154 520 158
rect 531 150 535 162
rect 542 154 550 158
rect 578 150 582 161
rect 589 154 596 158
rect -54 136 -33 141
rect -123 128 -103 132
rect -88 128 -79 132
rect -72 131 -61 132
rect -72 128 -56 131
rect -123 127 -119 128
rect -161 125 -157 126
rect -169 118 -165 121
rect -88 124 -84 128
rect -72 125 -68 128
rect -139 117 -135 119
rect -143 113 -135 117
rect -80 116 -76 121
rect -104 112 -100 116
rect -62 111 -56 128
rect -92 106 -88 109
rect -66 105 -56 111
rect -135 101 -131 104
rect -162 64 -158 67
rect -174 51 -170 60
rect -151 59 -135 63
rect -180 24 -173 28
rect -158 25 -154 35
rect -151 25 -147 59
rect -144 51 -140 56
rect -108 52 -105 56
rect -119 43 -115 52
rect -101 43 -97 49
rect -85 43 -81 49
rect -166 22 -147 25
rect -128 28 -124 35
rect -111 28 -107 35
rect -93 28 -89 35
rect -77 28 -73 35
rect -128 24 -108 28
rect -93 24 -84 28
rect -77 24 -69 28
rect -38 30 -33 136
rect -28 104 -23 148
rect 200 147 226 150
rect 247 147 265 150
rect 288 147 313 150
rect 328 147 347 150
rect 369 147 388 150
rect 409 147 430 150
rect 448 147 459 150
rect 490 147 510 150
rect 530 147 550 150
rect 571 147 591 150
rect -3 133 28 137
rect -3 132 1 133
rect -6 128 1 132
rect 24 129 31 133
rect 60 130 64 136
rect 307 134 313 147
rect 661 145 665 158
rect 679 157 691 161
rect 679 147 691 151
rect 643 143 665 145
rect 643 139 671 143
rect 700 143 704 158
rect 758 150 762 153
rect 332 134 338 137
rect 643 134 649 139
rect 26 126 29 129
rect 18 122 30 126
rect 107 128 649 134
rect 663 132 667 139
rect 682 138 686 140
rect 695 139 704 143
rect 700 133 704 139
rect 679 129 695 133
rect 699 129 704 133
rect 746 137 750 146
rect 769 145 785 149
rect 0 104 4 115
rect 18 114 30 118
rect 18 104 30 108
rect -28 100 4 104
rect -28 99 10 100
rect 0 96 10 99
rect 39 100 43 115
rect 55 108 60 114
rect 68 113 72 122
rect 307 113 313 128
rect 332 127 338 128
rect 663 121 671 125
rect 699 121 704 125
rect 68 108 483 113
rect 744 110 747 114
rect 762 111 766 121
rect 769 111 773 145
rect 776 137 780 142
rect 812 138 815 142
rect 801 129 805 138
rect 819 129 823 135
rect 835 129 839 135
rect 754 108 773 111
rect 792 114 796 121
rect 809 114 813 121
rect 827 114 831 121
rect 843 114 847 121
rect 792 110 812 114
rect 827 110 836 114
rect 843 110 854 114
rect 792 109 796 110
rect 68 105 72 108
rect 2 89 6 96
rect 21 95 25 97
rect 34 96 43 100
rect 60 96 64 101
rect 68 100 72 101
rect 68 96 77 100
rect 39 90 43 96
rect 18 86 34 90
rect 38 86 43 90
rect 2 78 10 82
rect 38 78 43 82
rect -9 58 29 65
rect 26 54 29 58
rect 60 58 64 64
rect 18 50 30 54
rect 307 55 313 108
rect 754 107 758 108
rect 746 100 750 103
rect 827 106 831 110
rect 843 107 847 110
rect 776 99 780 101
rect 772 95 780 99
rect 835 98 839 103
rect 811 94 815 98
rect 476 88 647 94
rect 641 60 647 88
rect 823 88 827 91
rect 696 82 699 86
rect 780 83 784 86
rect 688 78 700 82
rect 670 60 674 71
rect 688 70 700 74
rect 688 60 700 64
rect 641 56 674 60
rect 0 30 4 43
rect 18 42 30 46
rect 18 32 30 36
rect -38 28 4 30
rect -38 25 10 28
rect 0 24 10 25
rect 39 28 43 43
rect 68 42 72 50
rect 165 49 564 55
rect 641 54 680 56
rect 670 52 680 54
rect 709 56 713 71
rect 165 42 171 49
rect 55 36 60 42
rect 68 36 171 42
rect 68 33 72 36
rect -128 23 -124 24
rect -166 21 -162 22
rect -174 14 -170 17
rect -93 20 -89 24
rect -77 21 -73 24
rect -144 13 -140 15
rect -148 9 -140 13
rect 2 17 6 24
rect 21 23 25 25
rect 34 24 43 28
rect 60 24 64 29
rect 68 28 72 29
rect 68 24 77 28
rect 307 24 313 49
rect 672 45 676 52
rect 691 51 695 53
rect 704 52 713 56
rect 762 56 766 59
rect 709 46 713 52
rect 688 42 704 46
rect 708 42 713 46
rect 750 43 754 52
rect 773 51 789 55
rect 672 34 680 38
rect 708 34 713 38
rect 556 26 625 32
rect 39 18 43 24
rect -85 12 -81 17
rect 18 14 34 18
rect 38 14 43 18
rect -109 8 -105 12
rect 2 6 10 10
rect 38 6 43 10
rect -97 2 -93 5
rect -140 -3 -136 0
rect -168 -50 -164 -47
rect -180 -63 -176 -54
rect -157 -55 -141 -51
rect -186 -90 -179 -86
rect -164 -89 -160 -79
rect -157 -89 -153 -55
rect -150 -63 -146 -58
rect -114 -62 -111 -58
rect -125 -71 -121 -62
rect -107 -71 -103 -65
rect -91 -71 -87 -65
rect -172 -92 -153 -89
rect -134 -86 -130 -79
rect -117 -86 -113 -79
rect -99 -86 -95 -79
rect -83 -86 -79 -79
rect 619 -80 625 26
rect 747 16 751 20
rect 766 17 770 27
rect 773 17 777 51
rect 780 43 784 48
rect 816 44 819 48
rect 805 35 809 44
rect 823 35 827 41
rect 839 35 843 41
rect 758 14 777 17
rect 796 20 800 27
rect 813 20 817 27
rect 831 20 835 27
rect 847 20 851 27
rect 796 16 816 20
rect 831 16 840 20
rect 847 16 858 20
rect 796 15 800 16
rect 758 13 762 14
rect 750 6 754 9
rect 831 12 835 16
rect 847 13 851 16
rect 780 5 784 7
rect 776 1 784 5
rect 839 4 843 9
rect 815 0 819 4
rect 827 -6 831 -3
rect 784 -11 788 -8
rect 763 -43 767 -40
rect 696 -54 699 -50
rect 688 -58 700 -54
rect 751 -56 755 -47
rect 774 -48 790 -44
rect 670 -80 674 -65
rect 688 -66 700 -62
rect 688 -76 700 -72
rect -134 -90 -114 -86
rect -99 -90 -90 -86
rect -83 -90 -76 -86
rect 619 -84 680 -80
rect 709 -80 713 -65
rect 619 -86 676 -84
rect 691 -85 695 -83
rect 704 -84 713 -80
rect 749 -83 752 -79
rect 767 -82 771 -72
rect 774 -82 778 -48
rect 781 -56 785 -51
rect 817 -55 820 -51
rect 806 -64 810 -55
rect 824 -64 828 -58
rect 840 -64 844 -58
rect -134 -91 -130 -90
rect -172 -93 -168 -92
rect -180 -100 -176 -97
rect -99 -94 -95 -90
rect -83 -93 -79 -90
rect -150 -101 -146 -99
rect -154 -105 -146 -101
rect -91 -102 -87 -97
rect -115 -106 -111 -102
rect -103 -112 -99 -109
rect 257 -108 261 -86
rect 271 -96 291 -93
rect 271 -100 275 -96
rect 287 -100 291 -96
rect 279 -108 283 -104
rect 257 -111 283 -108
rect 311 -108 315 -86
rect 325 -96 345 -93
rect 325 -100 329 -96
rect 341 -100 345 -96
rect 333 -108 337 -104
rect 311 -111 337 -108
rect 359 -108 363 -86
rect 373 -96 393 -93
rect 373 -100 377 -96
rect 389 -100 393 -96
rect 381 -108 385 -104
rect 359 -111 385 -108
rect 407 -108 411 -86
rect 421 -96 441 -93
rect 421 -100 425 -96
rect 437 -100 441 -96
rect 429 -108 433 -104
rect 407 -111 433 -108
rect 466 -108 470 -86
rect 672 -91 676 -86
rect 709 -90 713 -84
rect 759 -85 778 -82
rect 797 -79 801 -72
rect 814 -79 818 -72
rect 832 -79 836 -72
rect 848 -79 852 -72
rect 797 -83 817 -79
rect 832 -83 841 -79
rect 848 -83 859 -79
rect 797 -84 801 -83
rect 759 -86 763 -85
rect 480 -96 500 -93
rect 688 -94 704 -90
rect 708 -94 713 -90
rect 751 -93 755 -90
rect 832 -87 836 -83
rect 848 -86 852 -83
rect 781 -94 785 -92
rect 480 -100 484 -96
rect 496 -100 500 -96
rect 777 -98 785 -94
rect 840 -95 844 -90
rect 672 -102 680 -98
rect 708 -102 713 -98
rect 816 -99 820 -95
rect 488 -108 492 -104
rect 466 -111 492 -108
rect 828 -105 832 -102
rect 785 -110 789 -107
rect 257 -112 275 -111
rect 311 -112 329 -111
rect 359 -112 377 -111
rect 407 -112 425 -111
rect 466 -112 484 -111
rect -146 -117 -142 -114
rect 271 -120 275 -112
rect 325 -120 329 -112
rect 373 -120 377 -112
rect 421 -120 425 -112
rect 480 -120 484 -112
rect 287 -144 291 -136
rect 341 -144 345 -136
rect 389 -144 393 -136
rect 437 -144 441 -136
rect 496 -144 500 -136
rect 275 -154 279 -151
rect 283 -154 287 -151
rect 329 -154 333 -151
rect 337 -154 341 -151
rect 377 -154 381 -151
rect 385 -154 389 -151
rect 425 -154 429 -151
rect 433 -154 437 -151
rect 484 -154 488 -151
rect 492 -154 496 -151
rect 765 -148 769 -145
rect 753 -161 757 -152
rect 776 -153 792 -149
rect -171 -183 -167 -180
rect -183 -196 -179 -187
rect -160 -188 -144 -184
rect -189 -223 -182 -219
rect -167 -222 -163 -212
rect -160 -222 -156 -188
rect 700 -184 749 -183
rect 700 -188 754 -184
rect 769 -187 773 -177
rect 776 -187 780 -153
rect 783 -161 787 -156
rect 819 -160 822 -156
rect 808 -169 812 -160
rect 826 -169 830 -163
rect 842 -169 846 -163
rect 700 -189 710 -188
rect 761 -190 780 -187
rect 799 -184 803 -177
rect 816 -184 820 -177
rect 834 -184 838 -177
rect 850 -184 854 -177
rect 799 -188 819 -184
rect 834 -188 843 -184
rect 850 -188 861 -184
rect 799 -189 803 -188
rect 761 -191 765 -190
rect -153 -196 -149 -191
rect -117 -195 -114 -191
rect -128 -204 -124 -195
rect 753 -198 757 -195
rect 834 -192 838 -188
rect 850 -191 854 -188
rect -110 -204 -106 -198
rect -94 -204 -90 -198
rect 783 -199 787 -197
rect 779 -203 787 -199
rect 842 -200 846 -195
rect 818 -204 822 -200
rect -175 -225 -156 -222
rect -137 -219 -133 -212
rect -120 -219 -116 -212
rect -102 -219 -98 -212
rect -86 -219 -82 -212
rect 830 -210 834 -207
rect 787 -215 791 -212
rect -79 -219 -36 -217
rect -137 -223 -117 -219
rect -102 -223 -93 -219
rect -86 -223 -36 -219
rect -137 -224 -133 -223
rect -175 -226 -171 -225
rect -183 -233 -179 -230
rect -102 -227 -98 -223
rect -86 -226 -82 -223
rect -79 -224 -36 -223
rect -153 -234 -149 -232
rect -157 -238 -149 -234
rect -94 -235 -90 -230
rect -118 -239 -114 -235
rect -106 -245 -102 -242
rect -149 -250 -145 -247
rect -172 -295 -168 -292
rect -184 -308 -180 -299
rect -161 -300 -145 -296
rect -190 -335 -183 -331
rect -168 -334 -164 -324
rect -161 -334 -157 -300
rect -154 -308 -150 -303
rect -118 -307 -115 -303
rect -129 -316 -125 -307
rect -111 -316 -107 -310
rect -95 -316 -91 -310
rect -176 -337 -157 -334
rect -138 -331 -134 -324
rect -121 -331 -117 -324
rect -103 -331 -99 -324
rect -87 -331 -83 -324
rect -71 -331 -67 -329
rect -138 -335 -118 -331
rect -103 -335 -94 -331
rect -87 -335 -67 -331
rect -138 -336 -134 -335
rect -176 -338 -172 -337
rect -184 -345 -180 -342
rect -103 -339 -99 -335
rect -87 -338 -83 -335
rect -71 -336 -67 -335
rect -154 -346 -150 -344
rect -158 -350 -150 -346
rect -95 -347 -91 -342
rect -119 -351 -115 -347
rect -107 -357 -103 -354
rect -150 -362 -146 -359
<< m2contact >>
rect 144 387 150 393
rect 224 386 231 393
rect 246 347 252 354
rect 25 331 32 338
rect 22 313 28 319
rect 51 313 57 319
rect 96 326 102 332
rect 19 272 26 279
rect 21 245 27 251
rect 46 245 53 251
rect 436 278 443 285
rect 313 246 318 251
rect 518 239 523 244
rect 1 200 8 207
rect 21 178 27 184
rect 47 178 54 184
rect 231 193 237 199
rect 275 194 280 199
rect 313 194 318 199
rect 196 168 202 174
rect 355 193 361 199
rect 437 193 442 199
rect 483 193 488 198
rect 518 193 523 199
rect 560 193 566 199
rect 682 311 688 317
rect 644 294 650 300
rect 738 301 744 307
rect 682 236 688 242
rect 629 218 635 224
rect 737 206 743 212
rect 231 153 237 159
rect 276 153 281 159
rect 311 153 317 159
rect 358 153 364 159
rect 389 153 395 159
rect 438 153 443 159
rect 597 168 603 174
rect 470 153 476 159
rect 520 153 525 159
rect 550 153 556 159
rect 596 153 601 159
rect -72 105 -66 111
rect -69 24 -62 31
rect -13 127 -6 134
rect 682 151 688 157
rect 101 128 107 134
rect 21 108 27 114
rect 48 108 55 114
rect 483 108 488 113
rect 738 110 744 116
rect -16 58 -9 65
rect 470 88 476 94
rect 691 64 697 70
rect 21 36 27 42
rect 564 49 570 55
rect 48 36 55 42
rect 550 26 556 32
rect 741 15 747 21
rect 691 -72 697 -66
rect -76 -90 -71 -85
rect 256 -86 262 -81
rect 310 -86 316 -81
rect 358 -86 364 -81
rect 406 -86 412 -81
rect 465 -86 471 -81
rect 743 -83 749 -78
rect 694 -189 700 -183
rect -36 -224 -29 -217
rect -67 -336 -60 -329
<< metal2 >>
rect 144 385 150 387
rect 144 380 145 385
rect 144 379 150 380
rect 224 365 231 386
rect 224 359 361 365
rect 25 338 32 350
rect 252 348 280 353
rect 102 326 237 332
rect 28 313 51 319
rect 37 300 41 313
rect 51 294 57 313
rect 110 302 181 308
rect 110 294 116 302
rect 51 288 116 294
rect 175 300 181 302
rect -59 272 19 279
rect -72 103 -66 105
rect -67 98 -66 103
rect -72 97 -66 98
rect -59 31 -52 272
rect 27 245 46 251
rect 47 224 53 245
rect 47 218 131 224
rect -62 24 -52 31
rect -47 200 1 207
rect -47 50 -40 200
rect 27 178 47 184
rect 47 158 53 178
rect 47 152 107 158
rect 101 134 107 152
rect -36 127 -13 134
rect -47 -85 -42 50
rect -71 -90 -42 -85
rect -36 -217 -29 127
rect 27 108 48 114
rect 101 112 107 128
rect 131 126 137 218
rect 175 139 181 294
rect 231 199 237 326
rect 275 199 280 348
rect 313 199 318 246
rect 355 199 361 359
rect 688 311 730 317
rect 724 307 730 311
rect 724 301 738 307
rect 630 295 631 300
rect 636 295 644 300
rect 630 294 644 295
rect 437 199 442 278
rect 518 199 523 239
rect 688 236 725 242
rect 621 219 622 224
rect 627 219 629 224
rect 621 218 629 219
rect 719 212 725 236
rect 719 206 737 212
rect 566 193 570 198
rect 195 168 196 174
rect 231 139 237 153
rect 276 150 281 153
rect 175 133 237 139
rect 311 126 317 153
rect 358 150 364 153
rect 131 120 317 126
rect 389 112 395 153
rect 438 150 443 153
rect 48 81 54 108
rect 101 106 395 112
rect 470 94 476 153
rect 483 113 488 193
rect 520 151 525 153
rect 165 88 470 94
rect 165 81 171 88
rect 48 75 171 81
rect -16 -311 -9 58
rect 27 36 48 42
rect 48 17 54 36
rect 550 32 556 153
rect 564 55 570 193
rect 603 168 630 174
rect 596 152 601 153
rect 165 26 550 30
rect 165 24 556 26
rect 165 17 171 24
rect 48 11 171 17
rect 257 -81 261 -77
rect 311 -81 315 -77
rect 359 -81 363 -77
rect 407 -81 411 -77
rect 466 -81 470 -77
rect 624 -183 630 168
rect 688 151 727 157
rect 721 116 727 151
rect 721 110 738 116
rect 721 106 727 110
rect 697 64 727 70
rect 721 21 727 64
rect 721 15 741 21
rect 697 -72 733 -66
rect 726 -78 733 -72
rect 726 -83 743 -78
rect 726 -85 749 -83
rect 624 -189 694 -183
rect -67 -318 -9 -311
rect -67 -329 -60 -318
<< m3contact >>
rect 145 380 150 385
rect 25 350 32 355
rect 175 294 181 300
rect -72 98 -67 103
rect 131 218 137 224
rect 631 295 636 300
rect 622 219 627 224
rect 190 168 195 174
rect 275 145 282 150
rect 357 144 365 150
rect 437 144 444 150
rect 519 146 526 151
rect 595 147 602 152
rect 256 -77 262 -72
rect 310 -77 316 -72
rect 358 -77 364 -72
rect 406 -77 412 -72
rect 465 -77 471 -72
<< metal3 >>
rect 144 385 151 386
rect 144 380 145 385
rect 150 380 151 385
rect 144 379 151 380
rect 24 355 33 356
rect -53 350 25 355
rect 32 350 33 355
rect -53 349 33 350
rect -73 103 -66 104
rect -53 103 -47 349
rect 130 224 138 225
rect 137 218 138 224
rect 130 217 138 218
rect 144 174 150 379
rect 174 300 182 301
rect 630 300 637 301
rect 174 294 175 300
rect 181 295 631 300
rect 636 295 637 300
rect 181 294 637 295
rect 174 293 182 294
rect 621 224 628 225
rect 621 219 622 224
rect 627 219 628 224
rect 621 218 628 219
rect 189 174 196 175
rect 144 168 190 174
rect 195 168 196 174
rect 189 167 196 168
rect -73 98 -72 103
rect -67 98 -47 103
rect -73 97 -47 98
rect 276 2 281 145
rect 358 2 364 144
rect 257 -2 281 2
rect 311 -2 364 2
rect 257 -72 261 -2
rect 311 -72 315 -2
rect 438 -14 443 144
rect 359 -18 443 -14
rect 359 -72 363 -18
rect 520 -24 525 146
rect 407 -29 525 -24
rect 407 -72 411 -29
rect 596 -40 601 147
rect 466 -44 601 -40
rect 466 -72 470 -44
<< m4contact >>
rect 125 218 131 224
rect 615 218 621 224
<< metal4 >>
rect 131 218 615 224
<< labels >>
rlabel metal1 41 284 43 285 7 GND
rlabel metal1 4 284 6 285 3 VDD
rlabel metal1 40 216 42 217 7 GND
rlabel metal1 3 216 5 217 3 VDD
rlabel metal1 40 149 42 150 7 GND
rlabel metal1 3 149 5 150 3 VDD
rlabel metal1 40 79 42 80 7 GND
rlabel metal1 3 79 5 80 3 VDD
rlabel metal1 40 7 42 8 7 GND
rlabel metal1 3 7 5 8 3 VDD
rlabel metal1 3 302 4 303 3 A1
rlabel metal1 24 300 25 301 1 B1
rlabel m2contact 28 332 29 333 1 B1
rlabel metal1 2 234 3 235 3 A2
rlabel metal1 23 232 24 233 1 B2
rlabel metal1 27 264 28 265 1 B2
rlabel metal1 2 167 3 168 3 A3
rlabel metal1 23 165 24 166 1 B3
rlabel metal1 27 197 28 198 1 B3
rlabel metal1 2 97 3 98 3 A4
rlabel metal1 27 127 28 128 1 B4
rlabel metal1 23 95 24 96 1 B4
rlabel metal1 2 25 3 26 3 A5
rlabel metal1 23 23 24 24 1 B5
rlabel metal1 27 55 28 56 1 B5
rlabel metal1 61 234 62 236 1 GND
rlabel metal1 61 167 62 169 1 GND
rlabel metal1 61 97 62 99 1 GND
rlabel metal1 61 25 62 27 1 GND
rlabel metal1 62 270 63 271 1 VDD
rlabel metal1 62 203 63 204 1 VDD
rlabel metal1 62 133 63 134 1 VDD
rlabel metal1 62 61 63 62 1 VDD
rlabel metal1 66 334 67 335 1 VDD
rlabel metal1 66 298 67 300 1 GND
rlabel metal1 157 372 158 373 1 GND
rlabel metal1 201 372 202 373 1 GND
rlabel metal1 245 372 246 373 1 GND
rlabel metal1 289 372 290 373 1 GND
rlabel metal1 333 372 334 373 1 GND
rlabel metal1 160 428 161 429 5 B1
rlabel metal1 169 428 170 429 5 A1
rlabel metal1 204 428 205 429 5 B2
rlabel metal1 213 428 214 429 5 A2
rlabel metal1 248 428 249 429 5 B3
rlabel metal1 257 428 258 429 5 A3
rlabel metal1 301 428 302 429 5 A4
rlabel metal1 292 428 293 429 5 B4
rlabel metal1 336 428 337 429 5 B5
rlabel metal1 345 428 346 429 5 A5
rlabel metal1 228 195 229 196 1 P1b
rlabel metal1 227 155 228 156 1 P1
rlabel m2contact 275 196 276 197 1 G1b
rlabel metal1 274 171 275 172 1 C1
rlabel metal1 307 156 308 157 1 P2
rlabel metal1 309 196 310 197 1 P2b
rlabel metal1 355 156 356 157 1 D2
rlabel m2contact 356 196 357 197 1 G2b
rlabel metal1 357 171 358 172 1 C2
rlabel metal1 390 196 391 197 1 P3b
rlabel metal1 439 171 440 172 1 C3
rlabel m2contact 437 196 438 197 1 G3b
rlabel metal1 436 156 437 157 1 D3
rlabel m2contact 471 156 472 157 1 P4
rlabel metal1 471 196 472 197 1 P4b
rlabel metal1 519 171 520 172 1 C4
rlabel m2contact 518 196 519 197 1 G4b
rlabel metal1 517 156 518 157 1 D4
rlabel metal1 552 196 553 197 1 P5b
rlabel m2contact 552 156 553 157 1 P5
rlabel metal1 599 196 600 197 7 G5b
rlabel m2contact 598 171 599 172 7 C5
rlabel metal1 385 156 386 157 1 P3
rlabel metal1 164 417 165 418 1 VDD
rlabel metal1 208 417 209 418 1 VDD
rlabel metal1 252 417 253 418 1 VDD
rlabel metal1 296 417 297 418 1 VDD
rlabel metal1 340 417 341 418 1 VDD
rlabel metal1 258 148 259 149 1 GND
rlabel metal1 342 148 343 149 1 GND
rlabel metal1 426 148 427 149 1 GND
rlabel metal1 505 148 506 149 1 GND
rlabel metal1 586 148 587 149 1 GND
rlabel metal1 583 204 584 205 1 VDD
rlabel metal1 504 204 505 205 1 VDD
rlabel metal1 425 204 426 205 1 VDD
rlabel metal1 343 204 344 205 1 VDD
rlabel metal1 258 204 259 205 1 VDD
rlabel metal1 274 156 275 157 1 D1
rlabel metal1 594 155 595 156 1 D5
rlabel metal1 490 -95 491 -94 1 GND
rlabel metal1 498 -143 499 -142 1 VDD
rlabel metal1 431 -95 432 -94 1 GND
rlabel metal1 439 -143 440 -142 1 VDD
rlabel metal1 391 -143 392 -142 1 VDD
rlabel metal1 383 -95 384 -94 1 GND
rlabel metal1 335 -95 336 -94 1 GND
rlabel metal1 343 -143 344 -142 1 VDD
rlabel metal1 289 -143 290 -142 1 VDD
rlabel metal1 281 -95 282 -94 1 GND
rlabel metal1 276 -153 277 -152 1 B1
rlabel metal1 285 -153 286 -152 1 A1
rlabel metal1 330 -153 331 -152 1 B2
rlabel metal1 339 -153 340 -152 1 A2
rlabel metal1 378 -153 379 -152 1 B3
rlabel metal1 387 -153 388 -152 1 A3
rlabel metal1 426 -153 427 -152 1 B4
rlabel metal1 435 -153 436 -152 1 A4
rlabel metal1 485 -153 486 -152 1 B5
rlabel metal1 494 -153 495 -152 1 A5
rlabel metal1 701 122 703 123 7 GND
rlabel metal1 664 122 666 123 3 VDD
rlabel metal1 701 207 703 208 7 GND
rlabel metal1 664 207 666 208 3 VDD
rlabel metal1 701 282 703 283 7 GND
rlabel metal1 664 282 666 283 3 VDD
rlabel metal1 710 35 712 36 7 GND
rlabel metal1 673 35 675 36 3 VDD
rlabel metal1 710 -101 712 -100 7 GND
rlabel metal1 673 -101 675 -100 3 VDD
rlabel metal1 663 300 664 301 1 P1
rlabel metal1 663 225 664 226 1 P2
rlabel metal1 663 140 664 141 1 P3
rlabel metal1 672 53 673 54 1 P4
rlabel metal1 672 -83 673 -82 1 P5
rlabel metal1 684 298 685 299 1 Cin
rlabel metal1 688 330 689 331 1 Cin
rlabel metal2 694 313 696 314 1 S1
rlabel metal1 688 255 689 256 1 C1
rlabel metal1 684 223 685 224 1 C1
rlabel metal2 698 238 699 239 1 S2
rlabel metal2 697 152 698 153 1 S3
rlabel metal2 707 65 708 66 1 S4
rlabel metal2 707 -70 708 -69 1 S5
rlabel metal1 688 170 689 171 1 C2
rlabel metal1 684 138 685 139 1 C2
rlabel metal1 697 83 698 84 1 C3
rlabel metal1 693 51 694 52 1 C3
rlabel metal1 697 -53 698 -52 1 C4
rlabel metal1 693 -85 694 -84 1 C4
rlabel metal1 858 -186 859 -185 7 C5f
rlabel metal1 839 -186 840 -185 1 C5fb
rlabel metal1 851 112 852 113 1 S3f
rlabel metal1 856 -81 857 -80 7 S5f
rlabel metal1 837 -81 838 -80 1 S5fb
rlabel metal1 855 18 856 19 1 S4f
rlabel metal1 836 18 837 19 1 S4fb
rlabel metal1 832 111 833 112 1 S3fb
rlabel metal1 850 208 851 209 1 S2f
rlabel metal1 831 208 832 209 1 S2fb
rlabel m2contact 746 17 747 18 1 S4
rlabel m2contact 741 206 742 207 1 S2
rlabel metal1 850 302 851 303 1 S1f
rlabel metal1 831 303 832 304 1 S1fb
rlabel metal1 754 -197 755 -196 1 gnd
rlabel metal1 754 -154 755 -153 1 Vdd
rlabel metal1 766 -147 767 -146 5 Clk
rlabel metal1 843 -199 844 -198 1 gnd
rlabel metal1 843 -165 844 -164 1 Vdd
rlabel metal1 819 -203 820 -202 1 gnd
rlabel metal1 828 -165 829 -164 1 Vdd
rlabel metal1 831 -209 832 -208 1 Clk
rlabel metal1 809 -162 810 -161 1 Vdd
rlabel metal1 820 -158 821 -157 1 Reset
rlabel metal1 784 -159 785 -158 1 Vdd
rlabel metal1 781 -202 782 -201 1 gnd
rlabel metal1 788 -214 789 -213 1 Clk
rlabel metal1 746 292 747 293 1 gnd
rlabel metal1 746 335 747 336 1 Vdd
rlabel metal1 758 342 759 343 5 Clk
rlabel metal1 835 290 836 291 1 gnd
rlabel metal1 835 324 836 325 1 Vdd
rlabel metal1 811 286 812 287 1 gnd
rlabel metal1 820 324 821 325 1 Vdd
rlabel metal1 823 280 824 281 1 Clk
rlabel metal1 801 327 802 328 1 Vdd
rlabel metal1 812 331 813 332 1 Reset
rlabel metal1 776 330 777 331 1 Vdd
rlabel metal1 773 287 774 288 1 gnd
rlabel metal1 780 275 781 276 1 Clk
rlabel metal1 746 197 747 198 1 gnd
rlabel metal1 746 240 747 241 1 Vdd
rlabel metal1 758 247 759 248 5 Clk
rlabel metal1 835 195 836 196 1 gnd
rlabel metal1 835 229 836 230 1 Vdd
rlabel metal1 811 191 812 192 1 gnd
rlabel metal1 820 229 821 230 1 Vdd
rlabel metal1 823 185 824 186 1 Clk
rlabel metal1 801 232 802 233 1 Vdd
rlabel metal1 812 236 813 237 1 Reset
rlabel metal1 776 235 777 236 1 Vdd
rlabel metal1 773 192 774 193 1 gnd
rlabel metal1 780 180 781 181 1 Clk
rlabel metal1 747 101 748 102 1 gnd
rlabel metal1 747 144 748 145 1 Vdd
rlabel metal1 759 151 760 152 5 Clk
rlabel metal1 836 99 837 100 1 gnd
rlabel metal1 836 133 837 134 1 Vdd
rlabel metal1 812 95 813 96 1 gnd
rlabel metal1 821 133 822 134 1 Vdd
rlabel metal1 824 89 825 90 1 Clk
rlabel metal1 802 136 803 137 1 Vdd
rlabel metal1 813 140 814 141 1 Reset
rlabel metal1 777 139 778 140 1 Vdd
rlabel metal1 774 96 775 97 1 gnd
rlabel metal1 781 84 782 85 1 Clk
rlabel metal1 785 -10 786 -9 1 Clk
rlabel metal1 778 2 779 3 1 gnd
rlabel metal1 781 45 782 46 1 Vdd
rlabel metal1 817 46 818 47 1 Reset
rlabel metal1 806 42 807 43 1 Vdd
rlabel metal1 828 -5 829 -4 1 Clk
rlabel metal1 825 39 826 40 1 Vdd
rlabel metal1 816 1 817 2 1 gnd
rlabel metal1 840 39 841 40 1 Vdd
rlabel metal1 840 5 841 6 1 gnd
rlabel metal1 763 57 764 58 5 Clk
rlabel metal1 751 50 752 51 1 Vdd
rlabel metal1 751 7 752 8 1 gnd
rlabel metal1 752 -92 753 -91 1 gnd
rlabel metal1 752 -49 753 -48 1 Vdd
rlabel metal1 764 -42 765 -41 5 Clk
rlabel metal1 841 -94 842 -93 1 gnd
rlabel metal1 841 -60 842 -59 1 Vdd
rlabel metal1 817 -98 818 -97 1 gnd
rlabel metal1 826 -60 827 -59 1 Vdd
rlabel metal1 829 -104 830 -103 1 Clk
rlabel metal1 807 -57 808 -56 1 Vdd
rlabel metal1 818 -53 819 -52 1 Reset
rlabel metal1 782 -54 783 -53 1 Vdd
rlabel metal1 779 -97 780 -96 1 gnd
rlabel metal1 786 -109 787 -108 1 Clk
rlabel m2contact 741 302 742 303 1 S1
rlabel m2contact 742 111 743 112 1 S3
rlabel m2contact 747 -82 748 -81 1 S5
rlabel metal1 749 -187 750 -186 1 C5
rlabel metal1 -94 -88 -93 -87 1 B3b
rlabel metal1 -88 26 -87 27 1 B2b
rlabel metal1 -83 130 -82 131 1 B1b
rlabel metal1 -64 130 -63 131 1 B1
rlabel m2contact -69 26 -68 27 1 B2
rlabel metal1 -184 -89 -183 -88 1 B3i
rlabel metal1 -178 25 -177 26 1 B2i
rlabel metal1 -173 129 -172 130 1 B1i
rlabel metal1 -145 -116 -144 -115 1 Clk
rlabel metal1 -152 -104 -151 -103 1 gnd
rlabel metal1 -149 -61 -148 -60 1 Vdd
rlabel metal1 -113 -60 -112 -59 1 Reset
rlabel metal1 -124 -64 -123 -63 1 Vdd
rlabel metal1 -102 -111 -101 -110 1 Clk
rlabel metal1 -105 -67 -104 -66 1 Vdd
rlabel metal1 -114 -105 -113 -104 1 gnd
rlabel metal1 -90 -67 -89 -66 1 Vdd
rlabel metal1 -90 -101 -89 -100 1 gnd
rlabel metal1 -167 -49 -166 -48 5 Clk
rlabel metal1 -179 -56 -178 -55 1 Vdd
rlabel metal1 -179 -99 -178 -98 1 gnd
rlabel metal1 -139 -2 -138 -1 1 Clk
rlabel metal1 -146 10 -145 11 1 gnd
rlabel metal1 -143 53 -142 54 1 Vdd
rlabel metal1 -107 54 -106 55 1 Reset
rlabel metal1 -118 50 -117 51 1 Vdd
rlabel metal1 -96 3 -95 4 1 Clk
rlabel metal1 -99 47 -98 48 1 Vdd
rlabel metal1 -108 9 -107 10 1 gnd
rlabel metal1 -84 47 -83 48 1 Vdd
rlabel metal1 -84 13 -83 14 1 gnd
rlabel metal1 -161 65 -160 66 5 Clk
rlabel metal1 -173 58 -172 59 1 Vdd
rlabel metal1 -173 15 -172 16 1 gnd
rlabel metal1 -168 119 -167 120 1 gnd
rlabel metal1 -168 162 -167 163 1 Vdd
rlabel metal1 -156 169 -155 170 5 Clk
rlabel metal1 -79 117 -78 118 1 gnd
rlabel metal1 -79 151 -78 152 1 Vdd
rlabel metal1 -103 113 -102 114 1 gnd
rlabel metal1 -94 151 -93 152 1 Vdd
rlabel metal1 -91 107 -90 108 1 Clk
rlabel metal1 -113 154 -112 155 1 Vdd
rlabel metal1 -102 158 -101 159 1 Reset
rlabel metal1 -138 157 -137 158 1 Vdd
rlabel metal1 -141 114 -140 115 1 gnd
rlabel metal1 -134 102 -133 103 1 Clk
rlabel metal1 -98 -333 -97 -332 1 B5b
rlabel metal1 -97 -221 -96 -220 1 B4b
rlabel metal1 -78 -221 -77 -220 1 B4
rlabel metal1 -188 -334 -187 -333 3 B5i
rlabel metal1 -187 -222 -186 -221 3 B4i
rlabel metal1 -149 -361 -148 -360 1 Clk
rlabel metal1 -156 -349 -155 -348 1 gnd
rlabel metal1 -153 -306 -152 -305 1 Vdd
rlabel metal1 -117 -305 -116 -304 1 Reset
rlabel metal1 -128 -309 -127 -308 1 Vdd
rlabel metal1 -106 -356 -105 -355 1 Clk
rlabel metal1 -109 -312 -108 -311 1 Vdd
rlabel metal1 -118 -350 -117 -349 1 gnd
rlabel metal1 -94 -312 -93 -311 1 Vdd
rlabel metal1 -94 -346 -93 -345 1 gnd
rlabel metal1 -171 -294 -170 -293 5 Clk
rlabel metal1 -183 -301 -182 -300 1 Vdd
rlabel metal1 -183 -344 -182 -343 1 gnd
rlabel metal1 -148 -249 -147 -248 1 Clk
rlabel metal1 -155 -237 -154 -236 1 gnd
rlabel metal1 -152 -194 -151 -193 1 Vdd
rlabel metal1 -116 -193 -115 -192 1 Reset
rlabel metal1 -127 -197 -126 -196 1 Vdd
rlabel metal1 -105 -244 -104 -243 1 Clk
rlabel metal1 -108 -200 -107 -199 1 Vdd
rlabel metal1 -117 -238 -116 -237 1 gnd
rlabel metal1 -93 -200 -92 -199 1 Vdd
rlabel metal1 -93 -234 -92 -233 1 gnd
rlabel metal1 -170 -182 -169 -181 5 Clk
rlabel metal1 -182 -189 -181 -188 1 Vdd
rlabel metal1 -182 -232 -181 -231 1 gnd
rlabel metal1 -84 206 -83 207 1 A5b
rlabel metal1 -85 305 -84 306 1 A4b
rlabel metal1 -89 398 -88 399 1 A3b
rlabel metal1 -90 590 -89 591 1 A1b
rlabel metal1 -90 495 -89 496 1 A2b
rlabel metal1 -71 589 -70 590 1 A1
rlabel metal1 -71 495 -70 496 1 A2
rlabel metal1 -70 399 -69 400 1 A3
rlabel metal1 -66 305 -65 306 1 A4
rlabel metal1 -65 206 -64 207 1 A5
rlabel metal1 -174 205 -173 206 1 A5i
rlabel metal1 -175 304 -174 305 1 A4i
rlabel metal1 -179 398 -178 399 1 A3i
rlabel metal1 -180 589 -179 590 1 A1i
rlabel metal1 -180 494 -179 495 1 A2i
rlabel metal1 -175 579 -174 580 1 gnd
rlabel metal1 -175 622 -174 623 1 Vdd
rlabel metal1 -163 629 -162 630 5 Clk
rlabel metal1 -86 577 -85 578 1 gnd
rlabel metal1 -86 611 -85 612 1 Vdd
rlabel metal1 -110 573 -109 574 1 gnd
rlabel metal1 -101 611 -100 612 1 Vdd
rlabel metal1 -98 567 -97 568 1 Clk
rlabel metal1 -120 614 -119 615 1 Vdd
rlabel metal1 -109 618 -108 619 1 Reset
rlabel metal1 -145 617 -144 618 1 Vdd
rlabel metal1 -148 574 -147 575 1 gnd
rlabel metal1 -141 562 -140 563 1 Clk
rlabel metal1 -175 484 -174 485 1 gnd
rlabel metal1 -175 527 -174 528 1 Vdd
rlabel metal1 -163 534 -162 535 5 Clk
rlabel metal1 -86 482 -85 483 1 gnd
rlabel metal1 -86 516 -85 517 1 Vdd
rlabel metal1 -110 478 -109 479 1 gnd
rlabel metal1 -101 516 -100 517 1 Vdd
rlabel metal1 -98 472 -97 473 1 Clk
rlabel metal1 -120 519 -119 520 1 Vdd
rlabel metal1 -109 523 -108 524 1 Reset
rlabel metal1 -145 522 -144 523 1 Vdd
rlabel metal1 -148 479 -147 480 1 gnd
rlabel metal1 -141 467 -140 468 1 Clk
rlabel metal1 -174 388 -173 389 1 gnd
rlabel metal1 -174 431 -173 432 1 Vdd
rlabel metal1 -162 438 -161 439 5 Clk
rlabel metal1 -85 386 -84 387 1 gnd
rlabel metal1 -85 420 -84 421 1 Vdd
rlabel metal1 -109 382 -108 383 1 gnd
rlabel metal1 -100 420 -99 421 1 Vdd
rlabel metal1 -97 376 -96 377 1 Clk
rlabel metal1 -119 423 -118 424 1 Vdd
rlabel metal1 -108 427 -107 428 1 Reset
rlabel metal1 -144 426 -143 427 1 Vdd
rlabel metal1 -147 383 -146 384 1 gnd
rlabel metal1 -140 371 -139 372 1 Clk
rlabel metal1 -136 277 -135 278 1 Clk
rlabel metal1 -143 289 -142 290 1 gnd
rlabel metal1 -140 332 -139 333 1 Vdd
rlabel metal1 -104 333 -103 334 1 Reset
rlabel metal1 -115 329 -114 330 1 Vdd
rlabel metal1 -93 282 -92 283 1 Clk
rlabel metal1 -96 326 -95 327 1 Vdd
rlabel metal1 -105 288 -104 289 1 gnd
rlabel metal1 -81 326 -80 327 1 Vdd
rlabel metal1 -81 292 -80 293 1 gnd
rlabel metal1 -158 344 -157 345 5 Clk
rlabel metal1 -170 337 -169 338 1 Vdd
rlabel metal1 -170 294 -169 295 1 gnd
rlabel metal1 -169 195 -168 196 1 gnd
rlabel metal1 -169 238 -168 239 1 Vdd
rlabel metal1 -157 245 -156 246 5 Clk
rlabel metal1 -80 193 -79 194 1 gnd
rlabel metal1 -80 227 -79 228 1 Vdd
rlabel metal1 -104 189 -103 190 1 gnd
rlabel metal1 -95 227 -94 228 1 Vdd
rlabel metal1 -92 183 -91 184 1 Clk
rlabel metal1 -114 230 -113 231 1 Vdd
rlabel metal1 -103 234 -102 235 1 Reset
rlabel metal1 -139 233 -138 234 1 Vdd
rlabel metal1 -142 190 -141 191 1 gnd
rlabel metal1 -135 178 -134 179 1 Clk
rlabel metal1 118 413 119 414 1 Cinb
rlabel metal1 28 412 29 413 1 Cini
rlabel metal1 137 412 138 413 1 Cin
rlabel metal1 33 402 34 403 1 gnd
rlabel metal1 33 445 34 446 1 Vdd
rlabel metal1 45 452 46 453 5 Clk
rlabel metal1 122 400 123 401 1 gnd
rlabel metal1 122 434 123 435 1 Vdd
rlabel metal1 98 396 99 397 1 gnd
rlabel metal1 107 434 108 435 1 Vdd
rlabel metal1 110 390 111 391 1 Clk
rlabel metal1 88 437 89 438 1 Vdd
rlabel metal1 99 441 100 442 1 Reset
rlabel metal1 63 440 64 441 1 Vdd
rlabel metal1 60 397 61 398 1 gnd
rlabel metal1 67 385 68 386 1 Clk
rlabel m2contact 199 170 200 171 3 Cin
rlabel metal1 -79 -333 -78 -332 1 B5
rlabel m2contact -75 -88 -74 -87 1 B3
<< end >>
