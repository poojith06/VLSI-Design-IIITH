* FO4 Inverter Chain Example (Measure Rise/Fall Times at C and D)
.include TSMC_180nm.txt
.param Wn=1.8u
.param Wp={2.5*Wn}
.param L=0.18u
.global gnd
.subckt inverter in out vdd gnd Wn={Wn} Wp={Wp} L={L}
M1 out in gnd gnd CMOSN W={Wn} L={L}
M2 out in vdd vdd CMOSP W={Wp} L={L}
.ends inverter
Vdd vdd gnd 1.8
Vin A gnd PWL(0n 0V 0.5n 1.8V 1.1n 1.8V 1.5n 0V 5n 0V)
Xinv1 A  B vdd gnd inverter Wn={Wn}        Wp={Wp}        L={L}
Xinv2 B  C vdd gnd inverter Wn={4*Wn}      Wp={4*Wp}      L={L}
Xinv3 C  D vdd gnd inverter Wn={16*Wn}     Wp={16*Wp}     L={L}
Xinv4 D  E vdd gnd inverter Wn={64*Wn}     Wp={64*Wp}     L={L}
Xinv5 E  F vdd gnd inverter Wn={256*Wn}    Wp={256*Wp}    L={L}
Cload F gnd 1p
.control
tran 10p 5n
set curplottitle="mididoddisaipoojith-2025122010-4-B"
plot v(C) v(D)
meas tran trC TRIG v(C) VAL=0.18 RISE=1 TARG v(C) VAL=1.62 RISE=1
meas tran tfC TRIG v(C) VAL=1.62 FALL=1 TARG v(C) VAL=0.18 FALL=1
meas tran trD TRIG v(D) VAL=0.18 RISE=1 TARG v(D) VAL=1.62 RISE=1
meas tran tfD TRIG v(D) VAL=1.62 FALL=1 TARG v(D) VAL=0.18 FALL=1
print trC tfC trD tfD
.endc
.end