magic
tech scmos
timestamp 1763216542
<< nwell >>
rect 10 20 72 28
rect 10 0 123 20
<< ntransistor >>
rect 21 -12 23 -8
rect 51 -14 53 -6
rect 59 -14 61 -6
rect 86 -17 88 -9
rect 94 -17 96 -9
rect 110 -12 112 -8
<< ptransistor >>
rect 21 6 23 22
rect 29 6 31 22
rect 51 6 53 22
rect 59 6 61 22
rect 76 6 78 14
rect 94 6 96 14
rect 110 6 112 14
<< ndiffusion >>
rect 20 -12 21 -8
rect 23 -12 24 -8
rect 50 -14 51 -6
rect 53 -14 54 -6
rect 58 -14 59 -6
rect 61 -14 62 -6
rect 85 -17 86 -9
rect 88 -17 89 -9
rect 93 -17 94 -9
rect 96 -17 97 -9
rect 109 -12 110 -8
rect 112 -12 113 -8
<< pdiffusion >>
rect 20 6 21 22
rect 23 6 24 22
rect 28 6 29 22
rect 31 6 32 22
rect 50 6 51 22
rect 53 6 54 22
rect 58 6 59 22
rect 61 6 62 22
rect 75 6 76 14
rect 78 6 79 14
rect 93 6 94 14
rect 96 6 97 14
rect 109 6 110 14
rect 112 6 113 14
<< ndcontact >>
rect 16 -12 20 -8
rect 24 -12 28 -8
rect 46 -14 50 -6
rect 54 -14 58 -6
rect 62 -14 66 -6
rect 81 -17 85 -9
rect 89 -17 93 -9
rect 97 -17 101 -9
rect 105 -12 109 -8
rect 113 -12 117 -8
<< pdcontact >>
rect 16 6 20 22
rect 24 6 28 22
rect 32 6 36 22
rect 46 6 50 22
rect 54 6 58 22
rect 62 6 66 22
rect 71 6 75 14
rect 79 6 83 14
rect 89 6 93 14
rect 97 6 101 14
rect 105 6 109 14
rect 113 6 117 14
<< polysilicon >>
rect 21 22 23 25
rect 29 22 31 31
rect 51 22 53 25
rect 59 22 61 34
rect 76 14 78 27
rect 94 14 96 20
rect 110 14 112 20
rect 21 -8 23 6
rect 29 -2 31 6
rect 51 -6 53 6
rect 59 -6 61 6
rect 76 0 78 6
rect 94 -1 96 6
rect 86 -3 96 -1
rect 21 -15 23 -12
rect 86 -9 88 -3
rect 94 -9 96 -6
rect 110 -8 112 6
rect 51 -25 53 -14
rect 59 -17 61 -14
rect 110 -16 112 -12
rect 86 -20 88 -17
rect 94 -20 96 -17
<< polycontact >>
rect 28 31 32 35
rect 55 30 59 34
rect 78 23 82 27
rect 17 -5 21 -1
rect 82 -5 86 -1
rect 106 -5 110 -1
rect 93 -24 97 -20
rect 50 -29 54 -25
<< metal1 >>
rect 28 35 32 38
rect 16 22 20 31
rect 39 30 55 34
rect 10 -5 17 -1
rect 32 -4 36 6
rect 39 -4 43 30
rect 46 22 50 27
rect 82 23 85 27
rect 71 14 75 23
rect 89 14 93 20
rect 105 14 109 20
rect 24 -7 43 -4
rect 62 -1 66 6
rect 79 -1 83 6
rect 97 -1 101 6
rect 113 -1 117 6
rect 62 -5 82 -1
rect 97 -5 106 -1
rect 113 -5 124 -1
rect 62 -6 66 -5
rect 24 -8 28 -7
rect 16 -15 20 -12
rect 97 -9 101 -5
rect 113 -8 117 -5
rect 46 -16 50 -14
rect 42 -20 50 -16
rect 105 -17 109 -12
rect 81 -21 85 -17
rect 93 -27 97 -24
rect 50 -32 54 -29
<< labels >>
rlabel metal1 51 -31 52 -30 1 Clk
rlabel metal1 44 -19 45 -18 1 gnd
rlabel metal1 47 24 48 25 1 Vdd
rlabel metal1 65 -3 66 -2 1 B
rlabel metal1 83 25 84 26 1 Reset
rlabel metal1 72 21 73 22 1 Vdd
rlabel metal1 94 -26 95 -25 1 Clk
rlabel metal1 91 18 92 19 1 Vdd
rlabel metal1 82 -20 83 -19 1 gnd
rlabel metal1 121 -3 122 -2 7 Q
rlabel metal1 106 18 107 19 1 Vdd
rlabel metal1 106 -16 107 -15 1 gnd
rlabel metal1 29 36 30 37 5 Clk
rlabel metal1 12 -4 13 -3 3 D
rlabel metal1 41 -6 42 -5 1 A
rlabel metal1 17 29 18 30 1 Vdd
rlabel metal1 17 -14 18 -13 1 gnd
rlabel metal1 102 -3 103 -2 1 Qb
<< end >>
