* FO4 Inverter Chain (measure propagation delays for I3 and I4)
.include TSMC_180nm.txt
.param Wn=1.8u
.param Wp={2.5*Wn}
.param L=0.18u
.subckt inverter in out vdd gnd Wn={Wn} Wp={Wp} L={L}
M1 out in gnd gnd CMOSN W={Wn} L={L}
M2 out in vdd vdd CMOSP W={Wp} L={L}
.ends inverter
Vdd vdd 0 1.8
Vin A 0 PWL(0n 0V 0.5n 1.8V 1.1n 1.8V 1.5n 0V 5n 0V)
Xinv1 A  B vdd 0 inverter Wn={Wn}        Wp={Wp}        L={L}
Xinv2 B  C vdd 0 inverter Wn={4*Wn}      Wp={4*Wp}      L={L}
Xinv3 C  D vdd 0 inverter Wn={16*Wn}     Wp={16*Wp}     L={L}
Xinv4 D  E vdd 0 inverter Wn={64*Wn}     Wp={64*Wp}     L={L}
Xinv5 E  F vdd 0 inverter Wn={256*Wn}    Wp={256*Wp}    L={L}
Cload F 0 1p
.control
tran 10p 5n
plot v(C) v(D)
meas tran tplh_i3 TRIG v(C) VAL=0.9 RISE=1 TARG v(D) VAL=0.9 RISE=1
meas tran tphl_i3 TRIG v(C) VAL=0.9 FALL=1 TARG v(D) VAL=0.9 FALL=1
meas tran tplh_i4 TRIG v(D) VAL=0.9 RISE=1 TARG v(E) VAL=0.9 RISE=1
meas tran tphl_i4 TRIG v(D) VAL=0.9 FALL=1 TARG v(E) VAL=0.9 FALL=1
let tpd_i3 =(tplh_i3 + tphl_i3)/2
let tpd_i4 =(tplh_i4 + tphl_i4)/2
print tpd_i3 tpd_i4
.endc
.end