magic
tech scmos
timestamp 1763182219
<< nwell >>
rect -7 -3 35 21
<< ntransistor >>
rect 4 -23 6 -15
rect 22 -23 24 -15
<< ptransistor >>
rect 4 5 6 13
rect 22 5 24 13
<< ndiffusion >>
rect 3 -23 4 -15
rect 6 -23 7 -15
rect 21 -23 22 -15
rect 24 -23 25 -15
<< pdiffusion >>
rect 3 5 4 13
rect 6 5 7 13
rect 21 5 22 13
rect 24 5 25 13
<< ndcontact >>
rect -1 -23 3 -15
rect 7 -23 11 -15
rect 17 -23 21 -15
rect 25 -23 29 -15
<< pdcontact >>
rect -1 5 3 13
rect 7 5 11 13
rect 17 5 21 13
rect 25 5 29 13
<< polysilicon >>
rect 4 13 6 17
rect 22 13 24 17
rect 4 -15 6 5
rect 22 -15 24 5
rect 4 -27 6 -23
rect 22 -27 24 -23
<< polycontact >>
rect 0 -10 4 -6
rect 18 -11 22 -7
<< metal1 >>
rect 8 23 12 31
rect -1 19 21 23
rect -1 13 3 19
rect 17 13 21 19
rect 7 0 11 5
rect 25 0 29 5
rect 7 -4 49 0
rect -11 -10 0 -6
rect 15 -11 18 -7
rect 25 -15 29 -4
rect -1 -36 3 -23
rect 7 -27 21 -23
<< labels >>
rlabel metal1 9 25 10 27 5 VDD
rlabel metal1 1 -33 2 -31 1 GND
rlabel metal1 40 -3 41 -1 1 OUT
rlabel metal1 -4 -9 -3 -7 1 IN1
rlabel metal1 16 -11 17 -9 1 IN2
<< end >>
