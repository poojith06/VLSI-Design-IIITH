* ==========================================================
*  5-stage Manchester Carry Chain - Pre-layout
* ==========================================================

.include TSMC_180nm.txt
VDD Vdd 0 1.8

V_Cin  Cin  0 1.8

V_P1   P1   0 1.8
V_P2   P2   0 1.8
V_P3   P3   0 1.8
V_P4   P4   0 1.8
V_P5   P5   0 1.8

V_P1b  P1b  0 0
V_P2b  P2b  0 0
V_P3b  P3b  0 0
V_P4b  P4b  0 0
V_P5b  P5b  0 0

V_G1b  G1b  0 1.8
V_G2b  G2b  0 1.8
V_G3b  G3b  0 1.8
V_G4b  G4b  0 1.8
V_G5b  G5b  0 1.8

V_D1   D1   0 0
V_D2   D2   0 0
V_D3   D3   0 0
V_D4   D4   0 0
V_D5   D5   0 0

* ==========================================================
* Stage 1
* ==========================================================
MpassN1 C1 P1 Cin 0 CMOSN W=0.36u L=0.18u
MpassP1 C1 P1b Cin Vdd CMOSP W=0.72u L=0.18u
Mp1     C1    G1b Vdd Vdd CMOSP W=0.72u L=0.18u
Mn1     C1    D1  0   0   CMOSN W=0.36u L=0.18u

* ==========================================================
* Stage 2
* ==========================================================
MpassN2 C2 P2 C1 0 CMOSN W=0.36u L=0.18u
MpassP2 C2 P2b C1 Vdd CMOSP W=0.72u L=0.18u
Mp2     C2    G2b Vdd Vdd CMOSP W=0.72u L=0.18u
Mn2     C2    D2  0   0   CMOSN W=0.36u L=0.18u

* ==========================================================
* Stage 3
* ==========================================================
MpassN3 C3 P3 C2 0 CMOSN W=0.36u L=0.18u
MpassP3 C3 P3b C2 Vdd CMOSP W=0.72u L=0.18u
Mp3     C3    G3b Vdd Vdd CMOSP W=0.72u L=0.18u
Mn3     C3    D3  0   0   CMOSN W=0.36u L=0.18u

* ==========================================================
* Stage 4
* ==========================================================
MpassN4 C4 P4 C3 0 CMOSN W=0.36u L=0.18u
MpassP4 C4 P4b C3 Vdd CMOSP W=0.72u L=0.18u
Mp4     C4    G4b Vdd Vdd CMOSP W=0.72u L=0.18u
Mn4     C4    D4  0   0   CMOSN W=0.36u L=0.18u

* ==========================================================
* Stage 5
* ==========================================================
MpassN5 C5 P5 C4 0 CMOSN W=0.36u L=0.18u
MpassP5 C5 P5b C4 Vdd CMOSP W=0.72u L=0.18u
Mp5     C5    G5b Vdd Vdd CMOSP W=0.72u L=0.18u
Mn5     C5    D5  0   0   CMOSN W=0.36u L=0.18u

.tran 1n 200n
.control
run
plot v(Cin) v(C1) v(C2) v(C3) v(C4) v(C5)
.endc
.end
