.include TSMC_180nm.txt
.param LAMBDA=0.09u
.param width_N={20*LAMBDA}

.global gnd

Vin vin gnd 1.8
VGS ctrl gnd 1.8

Cout vout gnd 10p 
.ic V(vout)=0

M1 vout ctrl vin gnd CMOSN W={width_N} L={2*LAMBDA} 
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
+ AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

.control
tran 1n 1u
plot V(vout) 
.endc
.end