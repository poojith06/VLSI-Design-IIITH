magic
tech scmos
timestamp 1725253593
<< nwell >>
rect -2 -3 22 16
<< ntransistor >>
rect 9 -18 11 -11
<< ptransistor >>
rect 9 3 11 10
<< ndiffusion >>
rect 8 -18 9 -11
rect 11 -18 12 -11
<< pdiffusion >>
rect 8 3 9 10
rect 11 3 12 10
<< ndcontact >>
rect 4 -18 8 -11
rect 12 -18 16 -11
<< pdcontact >>
rect 4 3 8 10
rect 12 3 16 10
<< polysilicon >>
rect 9 10 11 16
rect 9 -11 11 3
rect 9 -22 11 -18
<< polycontact >>
rect 5 -7 9 -3
<< metal1 >>
rect -2 16 22 23
rect 4 10 8 16
rect -8 -7 5 -3
rect 12 -11 16 3
rect 4 -23 8 -18
rect -2 -30 22 -23
<< labels >>
rlabel metal1 -7 -5 -7 -5 3 in
rlabel metal1 3 -30 9 -24 1 gnd
rlabel metal1 12 -7 16 -4 1 out
rlabel metal1 0 17 6 23 5 vdd
<< end >>
