.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd

Vdd	vdd	gnd	1.8
vclk clk gnd pulse 0 1.8 0ns 0ns 0ns 10ns 20ns
vin d gnd pulse 0 1.8 7ns 0ns 0ns 43ns 86ns
vrst rst gnd pulse 0 1.8 0ns 0ns 0ns 40ns 80ns

M1_P2 temp1 d vdd vdd  CMOSP   W={1.44u} L={0.18u}
M2_P1 A clk temp1 vdd  CMOSP   W={1.44u} L={0.18u}
M3_N1 A d gnd gnd  CMOSN   W={0.36u} L={0.18u}
M4_P3 temp2 clk vdd vdd  CMOSP   W={1.44u} L={0.18u}
M5_P7 B A temp2 vdd  CMOSP   W={1.44u} L={0.18u}
M6_N3 B A temp3 gnd  CMOSN   W={0.72u} L={0.18u}
M7_N2 temp3 clk gnd gnd  CMOSN   W={0.72u} L={0.18u}
M8_P4 B rst vdd vdd  CMOSP   W={0.72u} L={0.18u}
M9_P5 qb B vdd vdd  CMOSP   W={0.72u} L={0.18u}
M10_N5 qb clk temp4 gnd  CMOSN   W={0.72u} L={0.18u}
M11_N4 temp4 B gnd gnd  CMOSN   W={0.72u} L={0.18u}
M12_P6 q qb vdd vdd  CMOSP   W={0.72u} L={0.18u}
M13_N6 q qb gnd gnd  CMOSN   W={0.36u} L={0.18u}

.tran 0.1n 200n
.control
run
plot v(clk)+8  v(rst)+6 v(d)+4 v(q)+2 

.endc
.end




// .include TSMC_180nm.txt
// .param SUPPLY=1.8
// .param LAMBDA=0.09u
// .global gnd vdd

// * --- Power Supply ---
// Vdd vdd gnd 1.8

// * --- Stimulus (Inputs) ---
// * CLOCK: Period 20ns, Rises exactly at 10.0ns
// vclk clk gnd pulse 0 1.8 10ns 100ps 100ps 10ns 20ns

// * 2. DATA: Rises at 9.5ns
// * This means Data is ready 100ps before the Clock rises.
// vin d gnd pulse 0 1.8 9.5ns 100ps 100ps 20ns 40ns

// * RESET: Inactive (Logic 0)
// vrst rst gnd 0

// * --- MTSPC Circuit ---
// M1_P2 temp1 d vdd vdd   CMOSP   W={1.44u} L={0.18u}
// M2_P1 A clk temp1 vdd   CMOSP   W={1.44u} L={0.18u}
// M3_N1 A d gnd gnd       CMOSN   W={0.36u} L={0.18u}
// M4_P3 temp2 clk vdd vdd CMOSP   W={1.44u} L={0.18u}
// M5_P7 B A temp2 vdd     CMOSP   W={1.44u} L={0.18u}
// M6_N3 B A temp3 gnd     CMOSN   W={0.72u} L={0.18u}
// M7_N2 temp3 clk gnd gnd CMOSN   W={0.72u} L={0.18u}
// M8_P4 B rst vdd vdd     CMOSP   W={0.72u} L={0.18u}
// M9_P5 qb B vdd vdd      CMOSP   W={0.72u} L={0.18u}
// M10_N5 qb clk temp4 gnd CMOSN   W={0.72u} L={0.18u}
// M11_N4 temp4 B gnd gnd  CMOSN   W={0.72u} L={0.18u}
// M12_P6 q qb vdd vdd     CMOSP   W={0.72u} L={0.18u}
// M13_N6 q qb gnd gnd     CMOSN   W={0.36u} L={0.18u}

// * --- Simulation Setup ---
// .ic v(q)=0
// .ic v(qb)=1.8
// .tran 0.01n 20n

// .control
// run

// * --- Plotting ---
// * Plot D, Internal Node A, Clock, and Output Q
// plot v(d) v(a) v(clk) v(q)

// * --- MEASUREMENTS ---

// * 1. SETUP TIME (t_setup)
// * Measured as the delay from Data (Rising) to Internal Node A (Falling)
// * This represents the speed of the first stage.
// meas tran t_setup trig v(d) val=0.9 rise=1 targ v(a) val=0.9 fall=1

// * 2. CLOCK-TO-Q DELAY (Tpcq)
// * Measured from Clock (Rising) to Output Q (Rising)
// meas tran t_pcq trig v(clk) val=0.9 rise=1 targ v(q) val=0.9 rise=1

// echo " "
// echo "=========================================="
// echo " TIMING ANALYSIS RESULTS "
// echo "=========================================="
// print t_setup
// print t_pcq
// echo "=========================================="

// .endc
// .end




